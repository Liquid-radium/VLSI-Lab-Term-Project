* 2-to-4 Decoder Subcircuit
* Active-High outputs created inside

.include "t14y_tsmc_025_level3.txt"

.subckt DEC2to4 A B Y0 Y1 Y2 Y3 vdd gnd

*---------------- Power supply ----------------
Vdd vdd 0 5

*---------------- Input signals ----------------
Va a 0 PULSE(0 5 0 1n 1n 10n 20n)   ; A toggles faster
Vb b 0 PULSE(0 5 0 1n 1n 20n 40n)   ; B toggles slower

*---------------- Inverters for A and B bar ----------------
* A -> Abar
Mp1 Abar a vdd vdd CMOSP W=4u L=1u
Mn1 Abar a 0   0   CMOSN W=2u L=1u

* B -> Bbar
Mp2 Bbar b vdd vdd CMOSP W=4u L=1u
Mn2 Bbar b 0   0   CMOSN W=2u L=1u

*---------------- Decoder Outputs ----------------
* Y0 = Abar & Bbar
Mp3 Y0 Abar vdd vdd CMOSP W=4u L=1u
Mp4 Y0 Bbar vdd vdd CMOSP W=4u L=1u
Mn3 Y0 Abar n1 n1 CMOSN W=2u L=1u
Mn4 n1 Bbar 0   0   CMOSN W=2u L=1u

* Y1 = Abar & B
Mp5 Y1 Abar vdd vdd CMOSP W=4u L=1u
Mp6 Y1 b    vdd vdd CMOSP W=4u L=1u
Mn5 Y1 Abar n2 n2 CMOSN W=2u L=1u
Mn6 n2 b    0   0  CMOSN W=2u L=1u

* Y2 = A & Bbar
Mp7 Y2 a    vdd vdd CMOSP W=4u L=1u
Mp8 Y2 Bbar vdd vdd CMOSP W=4u L=1u
Mn7 Y2 a    n3 n3 CMOSN W=2u L=1u
Mn8 n3 Bbar 0   0  CMOSN W=2u L=1u

* Y3 = A & B
Mp9  Y3 a vdd vdd CMOSP W=4u L=1u
Mp10 Y3 b vdd vdd CMOSP W=4u L=1u
Mn9  Y3 a n4 n4 CMOSN W=2u L=1u
Mn10 n4 b 0   0 CMOSN W=2u L=1u

* --- Active-High Inverters for Decoder Outputs ---
* Y0h, Y1h, Y2h, Y3h are the new active-high wordlines
Myn0 Y0h Y0 0 0 CMOSN W=2u L=1u
Myp0 Y0h Y0 vdd vdd CMOSP W=4u L=1u

Myn1 Y1h Y1 0 0 CMOSN W=2u L=1u
Myp1 Y1h Y1 vdd vdd CMOSP W=4u L=1u

Myn2 Y2h Y2 0 0 CMOSN W=2u L=1u
Myp2 Y2h Y2 vdd vdd CMOSP W=4u L=1u

Myn3 Y3h Y3 0 0 CMOSN W=2u L=1u
Myp3 Y3h Y3 vdd vdd CMOSP W=4u L=1u

*---------------- Simulation control ----------------
.tran 1n 200n
.control
run
plot v(a) v(b) v(Y0) v(Y1) v(Y2) v(Y3)
.endc

.ends DEC2to4
