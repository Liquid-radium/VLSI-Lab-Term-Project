* 2-to-4 Decoder Subcircuit
* Active-High outputs created inside
.subckt DEC2to4 A B Y0 Y1 Y2 Y3 Y0h Y1h Y2h Y3h vdd gnd

*---------------- Inverters for A and B bar ----------------
Mp1 Abar a vdd vdd CMOSP W=4u L=1u
Mn1 Abar a gnd gnd CMOSN W=2u L=1u

Mp2 Bbar b vdd vdd CMOSP W=4u L=1u
Mn2 Bbar b gnd gnd CMOSN W=2u L=1u

*---------------- Decoder Outputs ----------------
* Y0 = Abar & Bbar
Mp3 Y0 Abar vdd vdd CMOSP W=4u L=1u
Mp4 Y0 Bbar vdd vdd CMOSP W=4u L=1u
Mn3 Y0 Abar n1 n1 CMOSN W=2u L=1u
Mn4 n1 Bbar gnd gnd CMOSN W=2u L=1u

* Y1 = Abar & B
Mp5 Y1 Abar vdd vdd CMOSP W=4u L=1u
Mp6 Y1 b    vdd vdd CMOSP W=4u L=1u
Mn5 Y1 Abar n2 n2 CMOSN W=2u L=1u
Mn6 n2 b    gnd gnd CMOSN W=2u L=1u

* Y2 = A & Bbar
Mp7 Y2 a    vdd vdd CMOSP W=4u L=1u
Mp8 Y2 Bbar vdd vdd CMOSP W=4u L=1u
Mn7 Y2 a    n3 n3 CMOSN W=2u L=1u
Mn8 n3 Bbar gnd gnd CMOSN W=2u L=1u

* Y3 = A & B
Mp9  Y3 a vdd vdd CMOSP W=4u L=1u
Mp10 Y3 b vdd vdd CMOSP W=4u L=1u
Mn9  Y3 a n4 n4 CMOSN W=2u L=1u
Mn10 n4 b gnd gnd CMOSN W=2u L=1u

* --- Active-High Inverters for Decoder Outputs ---
Myn0 Y0h Y0 gnd gnd CMOSN W=2u L=1u
Myp0 Y0h Y0 vdd vdd CMOSP W=4u L=1u

Myn1 Y1h Y1 gnd gnd CMOSN W=2u L=1u
Myp1 Y1h Y1 vdd vdd CMOSP W=4u L=1u

Myn2 Y2h Y2 gnd gnd CMOSN W=2u L=1u
Myp2 Y2h Y2 vdd vdd CMOSP W=4u L=1u

Myn3 Y3h Y3 gnd gnd CMOSN W=2u L=1u
Myp3 Y3h Y3 vdd vdd CMOSP W=4u L=1u

.ends DEC2to4
* End of decoder.cir