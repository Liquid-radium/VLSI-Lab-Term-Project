* 2-to-4 Decoder Subcircuit
* Active-High outputs created inside

.include "t14y_tsmc_025_level3.txt"

.subckt DEC2to4 A B Y0 Y1 Y2 Y3 vdd gnd

* --- Inverters ---
Mp1 Abar A vdd vdd CMOSP W=4u L=1u
Mn1 Abar A gnd gnd CMOSN W=2u L=1u
Mp2 Bbar B vdd vdd CMOSP W=4u L=1u
Mn2 Bbar B gnd gnd CMOSN W=2u L=1u

* --- NAND outputs (active-low) ---
Mp3 Y0 Abar vdd vdd CMOSP W=4u L=1u
Mp4 Y0 Bbar vdd vdd CMOSP W=4u L=1u
Mn3 Y0 Abar n1 n1 CMOSN W=2u L=1u
Mn4 n1 Bbar gnd gnd CMOSN W=2u L=1u

Mp5 Y1 Abar vdd vdd CMOSP W=4u L=1u
Mp6 Y1 B vdd vdd CMOSP W=4u L=1u
Mn5 Y1 Abar n2 n2 CMOSN W=2u L=1u
Mn6 n2 B gnd gnd CMOSN W=2u L=1u

Mp7 Y2 A vdd vdd CMOSP W=4u L=1u
Mp8 Y2 Bbar vdd vdd CMOSP W=4u L=1u
Mn7 Y2 A n3 n3 CMOSN W=2u L=1u
Mn8 n3 Bbar gnd gnd CMOSN W=2u L=1u

Mp9 Y3 A vdd vdd CMOSP W=4u L=1u
Mp10 Y3 B vdd vdd CMOSP W=4u L=1u
Mn9 Y3 A n4 n4 CMOSN W=2u L=1u
Mn10 n4 B gnd gnd CMOSN W=2u L=1u

* --- Active-High Outputs ---
Myn0 Y0h Y0 gnd gnd CMOSN W=2u L=1u
Myp0 Y0h Y0 vdd vdd CMOSP W=4u L=1u

Myn1 Y1h Y1 gnd gnd CMOSN W=2u L=1u
Myp1 Y1h Y1 vdd vdd CMOSP W=4u L=1u

Myn2 Y2h Y2 gnd gnd CMOSN W=2u L=1u
Myp2 Y2h Y2 vdd vdd CMOSP W=4u L=1u

Myn3 Y3h Y3 gnd gnd CMOSN W=2u L=1u
Myp3 Y3h Y3 vdd vdd CMOSP W=4u L=1u

.ends DEC2to4
