magic
tech scmos
timestamp 1760475277
<< ab >>
rect -131 3 -107 75
rect -69 5 -29 77
rect 5 5 85 77
rect 87 5 167 77
rect 168 5 248 77
rect 251 5 331 77
rect -131 -76 -107 -4
rect -68 -74 -28 -2
rect 5 -76 165 -4
rect 168 -76 328 -4
rect -67 -153 -27 -81
rect 5 -158 325 -86
rect -67 -235 -27 -163
rect 5 -236 325 -164
<< nwell >>
rect -136 35 -102 80
rect -74 37 -24 82
rect 0 37 336 82
rect -136 -81 -102 -36
rect -73 -76 -23 -34
rect -73 -79 -22 -76
rect -72 -121 -22 -79
rect -72 -240 -22 -195
rect 0 -81 333 -36
rect 0 -126 330 -81
rect 0 -241 330 -196
<< pwell >>
rect -136 -36 -102 35
rect -74 3 -24 37
rect -74 0 -23 3
rect -73 -34 -23 0
rect 0 1 336 37
rect 0 -36 333 1
rect -72 -195 -22 -121
rect 0 -196 330 -126
<< poly >>
rect 47 73 76 75
rect 40 65 42 70
rect 47 65 49 73
rect 57 65 59 69
rect 64 65 66 69
rect 74 65 76 73
rect 129 73 158 75
rect 122 65 124 70
rect 129 65 131 73
rect 139 65 141 69
rect 146 65 148 69
rect 156 65 158 73
rect 210 73 239 75
rect 203 65 205 70
rect 210 65 212 73
rect 220 65 222 69
rect 227 65 229 69
rect 237 65 239 73
rect 293 73 322 75
rect 286 65 288 70
rect 293 65 295 73
rect 303 65 305 69
rect 310 65 312 69
rect 320 65 322 73
rect -50 62 -44 64
rect -122 60 -116 62
rect -50 60 -48 62
rect -46 60 -44 62
rect -122 58 -120 60
rect -118 58 -116 60
rect -122 56 -116 58
rect -122 53 -120 56
rect -60 55 -58 60
rect -50 58 -44 60
rect -50 53 -48 58
rect -40 53 -38 58
rect 14 55 16 60
rect 24 55 26 60
rect 40 56 42 59
rect 36 54 42 56
rect 36 52 38 54
rect 40 52 42 54
rect 36 50 42 52
rect -122 29 -120 41
rect -60 40 -58 43
rect -50 40 -48 43
rect -60 38 -54 40
rect -60 36 -58 38
rect -56 36 -54 38
rect -50 37 -46 40
rect -60 34 -54 36
rect -60 26 -58 34
rect -122 18 -120 23
rect -48 23 -46 37
rect -40 32 -38 43
rect 14 40 16 43
rect 24 40 26 43
rect 14 38 36 40
rect -41 30 -35 32
rect -41 28 -39 30
rect -37 28 -35 30
rect -41 26 -35 28
rect -41 23 -39 26
rect -60 16 -58 20
rect 15 21 17 38
rect 29 36 32 38
rect 34 36 36 38
rect 29 34 36 36
rect 29 31 31 34
rect 40 25 42 50
rect 47 40 49 59
rect 96 55 98 60
rect 106 55 108 60
rect 122 56 124 59
rect 57 50 59 53
rect 53 48 59 50
rect 64 48 66 53
rect 53 46 55 48
rect 57 46 59 48
rect 53 44 59 46
rect 63 46 69 48
rect 63 44 65 46
rect 67 44 69 46
rect 63 42 69 44
rect 47 38 59 40
rect 46 32 52 34
rect 46 30 48 32
rect 50 30 52 32
rect 46 28 52 30
rect 47 25 49 28
rect 57 25 59 38
rect 64 25 66 42
rect 74 38 76 53
rect 118 54 124 56
rect 118 52 120 54
rect 122 52 124 54
rect 118 50 124 52
rect 96 40 98 43
rect 106 40 108 43
rect 96 38 118 40
rect 70 36 76 38
rect 70 34 72 36
rect 74 34 76 36
rect 70 32 76 34
rect 74 29 76 32
rect 29 20 31 25
rect -48 9 -46 14
rect -41 9 -39 14
rect 15 10 17 15
rect 40 14 42 19
rect 47 14 49 19
rect 57 14 59 19
rect 64 14 66 19
rect 74 18 76 23
rect 97 21 99 38
rect 111 36 114 38
rect 116 36 118 38
rect 111 34 118 36
rect 111 31 113 34
rect 122 25 124 50
rect 129 40 131 59
rect 177 55 179 60
rect 187 55 189 60
rect 203 56 205 59
rect 139 50 141 53
rect 135 48 141 50
rect 146 48 148 53
rect 135 46 137 48
rect 139 46 141 48
rect 135 44 141 46
rect 145 46 151 48
rect 145 44 147 46
rect 149 44 151 46
rect 145 42 151 44
rect 129 38 141 40
rect 128 32 134 34
rect 128 30 130 32
rect 132 30 134 32
rect 128 28 134 30
rect 129 25 131 28
rect 139 25 141 38
rect 146 25 148 42
rect 156 38 158 53
rect 199 54 205 56
rect 199 52 201 54
rect 203 52 205 54
rect 199 50 205 52
rect 177 40 179 43
rect 187 40 189 43
rect 177 38 199 40
rect 152 36 158 38
rect 152 34 154 36
rect 156 34 158 36
rect 152 32 158 34
rect 156 29 158 32
rect 111 20 113 25
rect 97 10 99 15
rect 122 14 124 19
rect 129 14 131 19
rect 139 14 141 19
rect 146 14 148 19
rect 156 18 158 23
rect 178 21 180 38
rect 192 36 195 38
rect 197 36 199 38
rect 192 34 199 36
rect 192 31 194 34
rect 203 25 205 50
rect 210 40 212 59
rect 260 55 262 60
rect 270 55 272 60
rect 286 56 288 59
rect 220 50 222 53
rect 216 48 222 50
rect 227 48 229 53
rect 216 46 218 48
rect 220 46 222 48
rect 216 44 222 46
rect 226 46 232 48
rect 226 44 228 46
rect 230 44 232 46
rect 226 42 232 44
rect 210 38 222 40
rect 209 32 215 34
rect 209 30 211 32
rect 213 30 215 32
rect 209 28 215 30
rect 210 25 212 28
rect 220 25 222 38
rect 227 25 229 42
rect 237 38 239 53
rect 282 54 288 56
rect 282 52 284 54
rect 286 52 288 54
rect 282 50 288 52
rect 260 40 262 43
rect 270 40 272 43
rect 260 38 282 40
rect 233 36 239 38
rect 233 34 235 36
rect 237 34 239 36
rect 233 32 239 34
rect 237 29 239 32
rect 192 20 194 25
rect 178 10 180 15
rect 203 14 205 19
rect 210 14 212 19
rect 220 14 222 19
rect 227 14 229 19
rect 237 18 239 23
rect 261 21 263 38
rect 275 36 278 38
rect 280 36 282 38
rect 275 34 282 36
rect 275 31 277 34
rect 286 25 288 50
rect 293 40 295 59
rect 303 50 305 53
rect 299 48 305 50
rect 310 48 312 53
rect 299 46 301 48
rect 303 46 305 48
rect 299 44 305 46
rect 309 46 315 48
rect 309 44 311 46
rect 313 44 315 46
rect 309 42 315 44
rect 293 38 305 40
rect 292 32 298 34
rect 292 30 294 32
rect 296 30 298 32
rect 292 28 298 30
rect 293 25 295 28
rect 303 25 305 38
rect 310 25 312 42
rect 320 38 322 53
rect 316 36 322 38
rect 316 34 318 36
rect 320 34 322 36
rect 316 32 322 34
rect 320 29 322 32
rect 275 20 277 25
rect 261 10 263 15
rect 286 14 288 19
rect 293 14 295 19
rect 303 14 305 19
rect 310 14 312 19
rect 320 18 322 23
rect -47 -11 -45 -6
rect -40 -11 -38 -6
rect -59 -17 -57 -13
rect -122 -24 -120 -19
rect 15 -14 17 -9
rect 40 -18 42 -13
rect 47 -18 49 -13
rect 57 -18 59 -13
rect 64 -18 66 -13
rect 95 -14 97 -9
rect -122 -42 -120 -30
rect -59 -31 -57 -23
rect -59 -33 -53 -31
rect -59 -35 -57 -33
rect -55 -35 -53 -33
rect -47 -34 -45 -20
rect -40 -23 -38 -20
rect -40 -25 -34 -23
rect -40 -27 -38 -25
rect -36 -27 -34 -25
rect -40 -29 -34 -27
rect -59 -37 -53 -35
rect -49 -37 -45 -34
rect -59 -40 -57 -37
rect -49 -40 -47 -37
rect -39 -40 -37 -29
rect 15 -37 17 -20
rect 29 -24 31 -19
rect 74 -22 76 -17
rect 120 -18 122 -13
rect 127 -18 129 -13
rect 137 -18 139 -13
rect 144 -18 146 -13
rect 178 -14 180 -9
rect 29 -33 31 -30
rect 29 -35 36 -33
rect 29 -37 32 -35
rect 34 -37 36 -35
rect 14 -39 36 -37
rect 14 -42 16 -39
rect 24 -42 26 -39
rect -122 -57 -120 -54
rect -59 -57 -57 -52
rect -49 -55 -47 -50
rect -39 -55 -37 -50
rect 40 -49 42 -24
rect 47 -27 49 -24
rect 46 -29 52 -27
rect 46 -31 48 -29
rect 50 -31 52 -29
rect 46 -33 52 -31
rect 57 -37 59 -24
rect 36 -51 42 -49
rect 36 -53 38 -51
rect 40 -53 42 -51
rect -49 -57 -43 -55
rect -122 -59 -116 -57
rect -122 -61 -120 -59
rect -118 -61 -116 -59
rect -49 -59 -47 -57
rect -45 -59 -43 -57
rect 14 -59 16 -54
rect 24 -59 26 -54
rect 36 -55 42 -53
rect 40 -58 42 -55
rect 47 -39 59 -37
rect 47 -58 49 -39
rect 64 -41 66 -24
rect 74 -31 76 -28
rect 70 -33 76 -31
rect 70 -35 72 -33
rect 74 -35 76 -33
rect 70 -37 76 -35
rect 95 -37 97 -20
rect 109 -24 111 -19
rect 154 -22 156 -17
rect 203 -18 205 -13
rect 210 -18 212 -13
rect 220 -18 222 -13
rect 227 -18 229 -13
rect 258 -14 260 -9
rect 109 -33 111 -30
rect 109 -35 116 -33
rect 109 -37 112 -35
rect 114 -37 116 -35
rect 63 -43 69 -41
rect 53 -45 59 -43
rect 53 -47 55 -45
rect 57 -47 59 -45
rect 63 -45 65 -43
rect 67 -45 69 -43
rect 63 -47 69 -45
rect 53 -49 59 -47
rect 57 -52 59 -49
rect 64 -52 66 -47
rect 74 -52 76 -37
rect 94 -39 116 -37
rect 94 -42 96 -39
rect 104 -42 106 -39
rect -49 -61 -43 -59
rect -122 -63 -116 -61
rect 120 -49 122 -24
rect 127 -27 129 -24
rect 126 -29 132 -27
rect 126 -31 128 -29
rect 130 -31 132 -29
rect 126 -33 132 -31
rect 137 -37 139 -24
rect 116 -51 122 -49
rect 116 -53 118 -51
rect 120 -53 122 -51
rect 94 -59 96 -54
rect 104 -59 106 -54
rect 116 -55 122 -53
rect 120 -58 122 -55
rect 127 -39 139 -37
rect 127 -58 129 -39
rect 144 -41 146 -24
rect 154 -31 156 -28
rect 150 -33 156 -31
rect 150 -35 152 -33
rect 154 -35 156 -33
rect 150 -37 156 -35
rect 178 -37 180 -20
rect 192 -24 194 -19
rect 237 -22 239 -17
rect 283 -18 285 -13
rect 290 -18 292 -13
rect 300 -18 302 -13
rect 307 -18 309 -13
rect 192 -33 194 -30
rect 192 -35 199 -33
rect 192 -37 195 -35
rect 197 -37 199 -35
rect 143 -43 149 -41
rect 133 -45 139 -43
rect 133 -47 135 -45
rect 137 -47 139 -45
rect 143 -45 145 -43
rect 147 -45 149 -43
rect 143 -47 149 -45
rect 133 -49 139 -47
rect 137 -52 139 -49
rect 144 -52 146 -47
rect 154 -52 156 -37
rect 177 -39 199 -37
rect 177 -42 179 -39
rect 187 -42 189 -39
rect 203 -49 205 -24
rect 210 -27 212 -24
rect 209 -29 215 -27
rect 209 -31 211 -29
rect 213 -31 215 -29
rect 209 -33 215 -31
rect 220 -37 222 -24
rect 199 -51 205 -49
rect 199 -53 201 -51
rect 203 -53 205 -51
rect 177 -59 179 -54
rect 187 -59 189 -54
rect 199 -55 205 -53
rect 203 -58 205 -55
rect 210 -39 222 -37
rect 210 -58 212 -39
rect 227 -41 229 -24
rect 237 -31 239 -28
rect 233 -33 239 -31
rect 233 -35 235 -33
rect 237 -35 239 -33
rect 233 -37 239 -35
rect 258 -37 260 -20
rect 272 -24 274 -19
rect 317 -22 319 -17
rect 272 -33 274 -30
rect 272 -35 279 -33
rect 272 -37 275 -35
rect 277 -37 279 -35
rect 226 -43 232 -41
rect 216 -45 222 -43
rect 216 -47 218 -45
rect 220 -47 222 -45
rect 226 -45 228 -43
rect 230 -45 232 -43
rect 226 -47 232 -45
rect 216 -49 222 -47
rect 220 -52 222 -49
rect 227 -52 229 -47
rect 237 -52 239 -37
rect 257 -39 279 -37
rect 257 -42 259 -39
rect 267 -42 269 -39
rect 283 -49 285 -24
rect 290 -27 292 -24
rect 289 -29 295 -27
rect 289 -31 291 -29
rect 293 -31 295 -29
rect 289 -33 295 -31
rect 300 -37 302 -24
rect 279 -51 285 -49
rect 279 -53 281 -51
rect 283 -53 285 -51
rect 257 -59 259 -54
rect 267 -59 269 -54
rect 279 -55 285 -53
rect 283 -58 285 -55
rect 290 -39 302 -37
rect 290 -58 292 -39
rect 307 -41 309 -24
rect 317 -31 319 -28
rect 313 -33 319 -31
rect 313 -35 315 -33
rect 317 -35 319 -33
rect 313 -37 319 -35
rect 306 -43 312 -41
rect 296 -45 302 -43
rect 296 -47 298 -45
rect 300 -47 302 -45
rect 306 -45 308 -43
rect 310 -45 312 -43
rect 306 -47 312 -45
rect 296 -49 302 -47
rect 300 -52 302 -49
rect 307 -52 309 -47
rect 317 -52 319 -37
rect 40 -69 42 -64
rect 47 -72 49 -64
rect 57 -68 59 -64
rect 64 -68 66 -64
rect 74 -72 76 -64
rect 47 -74 76 -72
rect 120 -69 122 -64
rect 127 -72 129 -64
rect 137 -68 139 -64
rect 144 -68 146 -64
rect 154 -72 156 -64
rect 127 -74 156 -72
rect 203 -69 205 -64
rect 210 -72 212 -64
rect 220 -68 222 -64
rect 227 -68 229 -64
rect 237 -72 239 -64
rect 210 -74 239 -72
rect 283 -69 285 -64
rect 290 -72 292 -64
rect 300 -68 302 -64
rect 307 -68 309 -64
rect 317 -72 319 -64
rect 290 -74 319 -72
rect 47 -90 76 -88
rect -48 -96 -42 -94
rect -48 -98 -46 -96
rect -44 -98 -42 -96
rect 40 -98 42 -93
rect 47 -98 49 -90
rect 57 -98 59 -94
rect 64 -98 66 -94
rect 74 -98 76 -90
rect 127 -90 156 -88
rect 120 -98 122 -93
rect 127 -98 129 -90
rect 137 -98 139 -94
rect 144 -98 146 -94
rect 154 -98 156 -90
rect 207 -90 236 -88
rect 200 -98 202 -93
rect 207 -98 209 -90
rect 217 -98 219 -94
rect 224 -98 226 -94
rect 234 -98 236 -90
rect 287 -90 316 -88
rect 280 -98 282 -93
rect 287 -98 289 -90
rect 297 -98 299 -94
rect 304 -98 306 -94
rect 314 -98 316 -90
rect -58 -103 -56 -98
rect -48 -100 -42 -98
rect -48 -105 -46 -100
rect -38 -105 -36 -100
rect 14 -108 16 -103
rect 24 -108 26 -103
rect 40 -107 42 -104
rect -58 -118 -56 -115
rect -48 -118 -46 -115
rect -58 -120 -52 -118
rect -58 -122 -56 -120
rect -54 -122 -52 -120
rect -48 -121 -44 -118
rect -58 -124 -52 -122
rect -58 -132 -56 -124
rect -46 -135 -44 -121
rect -38 -126 -36 -115
rect 36 -109 42 -107
rect 36 -111 38 -109
rect 40 -111 42 -109
rect 36 -113 42 -111
rect 14 -123 16 -120
rect 24 -123 26 -120
rect 14 -125 36 -123
rect -39 -128 -33 -126
rect -39 -130 -37 -128
rect -35 -130 -33 -128
rect -39 -132 -33 -130
rect -39 -135 -37 -132
rect -58 -142 -56 -138
rect 15 -142 17 -125
rect 29 -127 32 -125
rect 34 -127 36 -125
rect 29 -129 36 -127
rect 29 -132 31 -129
rect 40 -138 42 -113
rect 47 -123 49 -104
rect 94 -108 96 -103
rect 104 -108 106 -103
rect 120 -107 122 -104
rect 57 -113 59 -110
rect 53 -115 59 -113
rect 64 -115 66 -110
rect 53 -117 55 -115
rect 57 -117 59 -115
rect 53 -119 59 -117
rect 63 -117 69 -115
rect 63 -119 65 -117
rect 67 -119 69 -117
rect 63 -121 69 -119
rect 47 -125 59 -123
rect 46 -131 52 -129
rect 46 -133 48 -131
rect 50 -133 52 -131
rect 46 -135 52 -133
rect 47 -138 49 -135
rect 57 -138 59 -125
rect 64 -138 66 -121
rect 74 -125 76 -110
rect 116 -109 122 -107
rect 116 -111 118 -109
rect 120 -111 122 -109
rect 116 -113 122 -111
rect 94 -123 96 -120
rect 104 -123 106 -120
rect 94 -125 116 -123
rect 70 -127 76 -125
rect 70 -129 72 -127
rect 74 -129 76 -127
rect 70 -131 76 -129
rect 74 -134 76 -131
rect -46 -149 -44 -144
rect -39 -149 -37 -144
rect 29 -143 31 -138
rect 15 -153 17 -148
rect 40 -149 42 -144
rect 47 -149 49 -144
rect 57 -149 59 -144
rect 64 -149 66 -144
rect 74 -145 76 -140
rect 95 -142 97 -125
rect 109 -127 112 -125
rect 114 -127 116 -125
rect 109 -129 116 -127
rect 109 -132 111 -129
rect 120 -138 122 -113
rect 127 -123 129 -104
rect 174 -108 176 -103
rect 184 -108 186 -103
rect 200 -107 202 -104
rect 137 -113 139 -110
rect 133 -115 139 -113
rect 144 -115 146 -110
rect 133 -117 135 -115
rect 137 -117 139 -115
rect 133 -119 139 -117
rect 143 -117 149 -115
rect 143 -119 145 -117
rect 147 -119 149 -117
rect 143 -121 149 -119
rect 127 -125 139 -123
rect 126 -131 132 -129
rect 126 -133 128 -131
rect 130 -133 132 -131
rect 126 -135 132 -133
rect 127 -138 129 -135
rect 137 -138 139 -125
rect 144 -138 146 -121
rect 154 -125 156 -110
rect 196 -109 202 -107
rect 196 -111 198 -109
rect 200 -111 202 -109
rect 196 -113 202 -111
rect 174 -123 176 -120
rect 184 -123 186 -120
rect 174 -125 196 -123
rect 150 -127 156 -125
rect 150 -129 152 -127
rect 154 -129 156 -127
rect 150 -131 156 -129
rect 154 -134 156 -131
rect 109 -143 111 -138
rect 95 -153 97 -148
rect 120 -149 122 -144
rect 127 -149 129 -144
rect 137 -149 139 -144
rect 144 -149 146 -144
rect 154 -145 156 -140
rect 175 -142 177 -125
rect 189 -127 192 -125
rect 194 -127 196 -125
rect 189 -129 196 -127
rect 189 -132 191 -129
rect 200 -138 202 -113
rect 207 -123 209 -104
rect 254 -108 256 -103
rect 264 -108 266 -103
rect 280 -107 282 -104
rect 217 -113 219 -110
rect 213 -115 219 -113
rect 224 -115 226 -110
rect 213 -117 215 -115
rect 217 -117 219 -115
rect 213 -119 219 -117
rect 223 -117 229 -115
rect 223 -119 225 -117
rect 227 -119 229 -117
rect 223 -121 229 -119
rect 207 -125 219 -123
rect 206 -131 212 -129
rect 206 -133 208 -131
rect 210 -133 212 -131
rect 206 -135 212 -133
rect 207 -138 209 -135
rect 217 -138 219 -125
rect 224 -138 226 -121
rect 234 -125 236 -110
rect 276 -109 282 -107
rect 276 -111 278 -109
rect 280 -111 282 -109
rect 276 -113 282 -111
rect 254 -123 256 -120
rect 264 -123 266 -120
rect 254 -125 276 -123
rect 230 -127 236 -125
rect 230 -129 232 -127
rect 234 -129 236 -127
rect 230 -131 236 -129
rect 234 -134 236 -131
rect 189 -143 191 -138
rect 175 -153 177 -148
rect 200 -149 202 -144
rect 207 -149 209 -144
rect 217 -149 219 -144
rect 224 -149 226 -144
rect 234 -145 236 -140
rect 255 -142 257 -125
rect 269 -127 272 -125
rect 274 -127 276 -125
rect 269 -129 276 -127
rect 269 -132 271 -129
rect 280 -138 282 -113
rect 287 -123 289 -104
rect 297 -113 299 -110
rect 293 -115 299 -113
rect 304 -115 306 -110
rect 293 -117 295 -115
rect 297 -117 299 -115
rect 293 -119 299 -117
rect 303 -117 309 -115
rect 303 -119 305 -117
rect 307 -119 309 -117
rect 303 -121 309 -119
rect 287 -125 299 -123
rect 286 -131 292 -129
rect 286 -133 288 -131
rect 290 -133 292 -131
rect 286 -135 292 -133
rect 287 -138 289 -135
rect 297 -138 299 -125
rect 304 -138 306 -121
rect 314 -125 316 -110
rect 310 -127 316 -125
rect 310 -129 312 -127
rect 314 -129 316 -127
rect 310 -131 316 -129
rect 314 -134 316 -131
rect 269 -143 271 -138
rect 255 -153 257 -148
rect 280 -149 282 -144
rect 287 -149 289 -144
rect 297 -149 299 -144
rect 304 -149 306 -144
rect 314 -145 316 -140
rect -46 -172 -44 -167
rect -39 -172 -37 -167
rect -58 -178 -56 -174
rect 15 -174 17 -169
rect 40 -178 42 -173
rect 47 -178 49 -173
rect 57 -178 59 -173
rect 64 -178 66 -173
rect 95 -174 97 -169
rect -58 -192 -56 -184
rect -58 -194 -52 -192
rect -58 -196 -56 -194
rect -54 -196 -52 -194
rect -46 -195 -44 -181
rect -39 -184 -37 -181
rect -39 -186 -33 -184
rect -39 -188 -37 -186
rect -35 -188 -33 -186
rect -39 -190 -33 -188
rect -58 -198 -52 -196
rect -48 -198 -44 -195
rect -58 -201 -56 -198
rect -48 -201 -46 -198
rect -38 -201 -36 -190
rect 15 -197 17 -180
rect 29 -184 31 -179
rect 74 -182 76 -177
rect 120 -178 122 -173
rect 127 -178 129 -173
rect 137 -178 139 -173
rect 144 -178 146 -173
rect 175 -174 177 -169
rect 29 -193 31 -190
rect 29 -195 36 -193
rect 29 -197 32 -195
rect 34 -197 36 -195
rect 14 -199 36 -197
rect 14 -202 16 -199
rect 24 -202 26 -199
rect -58 -218 -56 -213
rect -48 -216 -46 -211
rect -38 -216 -36 -211
rect 40 -209 42 -184
rect 47 -187 49 -184
rect 46 -189 52 -187
rect 46 -191 48 -189
rect 50 -191 52 -189
rect 46 -193 52 -191
rect 57 -197 59 -184
rect 36 -211 42 -209
rect 36 -213 38 -211
rect 40 -213 42 -211
rect -48 -218 -42 -216
rect -48 -220 -46 -218
rect -44 -220 -42 -218
rect 14 -219 16 -214
rect 24 -219 26 -214
rect 36 -215 42 -213
rect 40 -218 42 -215
rect 47 -199 59 -197
rect 47 -218 49 -199
rect 64 -201 66 -184
rect 74 -191 76 -188
rect 70 -193 76 -191
rect 70 -195 72 -193
rect 74 -195 76 -193
rect 70 -197 76 -195
rect 95 -197 97 -180
rect 109 -184 111 -179
rect 154 -182 156 -177
rect 200 -178 202 -173
rect 207 -178 209 -173
rect 217 -178 219 -173
rect 224 -178 226 -173
rect 255 -174 257 -169
rect 109 -193 111 -190
rect 109 -195 116 -193
rect 109 -197 112 -195
rect 114 -197 116 -195
rect 63 -203 69 -201
rect 53 -205 59 -203
rect 53 -207 55 -205
rect 57 -207 59 -205
rect 63 -205 65 -203
rect 67 -205 69 -203
rect 63 -207 69 -205
rect 53 -209 59 -207
rect 57 -212 59 -209
rect 64 -212 66 -207
rect 74 -212 76 -197
rect 94 -199 116 -197
rect 94 -202 96 -199
rect 104 -202 106 -199
rect -48 -222 -42 -220
rect 120 -209 122 -184
rect 127 -187 129 -184
rect 126 -189 132 -187
rect 126 -191 128 -189
rect 130 -191 132 -189
rect 126 -193 132 -191
rect 137 -197 139 -184
rect 116 -211 122 -209
rect 116 -213 118 -211
rect 120 -213 122 -211
rect 94 -219 96 -214
rect 104 -219 106 -214
rect 116 -215 122 -213
rect 120 -218 122 -215
rect 127 -199 139 -197
rect 127 -218 129 -199
rect 144 -201 146 -184
rect 154 -191 156 -188
rect 150 -193 156 -191
rect 150 -195 152 -193
rect 154 -195 156 -193
rect 150 -197 156 -195
rect 175 -197 177 -180
rect 189 -184 191 -179
rect 234 -182 236 -177
rect 280 -178 282 -173
rect 287 -178 289 -173
rect 297 -178 299 -173
rect 304 -178 306 -173
rect 189 -193 191 -190
rect 189 -195 196 -193
rect 189 -197 192 -195
rect 194 -197 196 -195
rect 143 -203 149 -201
rect 133 -205 139 -203
rect 133 -207 135 -205
rect 137 -207 139 -205
rect 143 -205 145 -203
rect 147 -205 149 -203
rect 143 -207 149 -205
rect 133 -209 139 -207
rect 137 -212 139 -209
rect 144 -212 146 -207
rect 154 -212 156 -197
rect 174 -199 196 -197
rect 174 -202 176 -199
rect 184 -202 186 -199
rect 200 -209 202 -184
rect 207 -187 209 -184
rect 206 -189 212 -187
rect 206 -191 208 -189
rect 210 -191 212 -189
rect 206 -193 212 -191
rect 217 -197 219 -184
rect 196 -211 202 -209
rect 196 -213 198 -211
rect 200 -213 202 -211
rect 174 -219 176 -214
rect 184 -219 186 -214
rect 196 -215 202 -213
rect 200 -218 202 -215
rect 207 -199 219 -197
rect 207 -218 209 -199
rect 224 -201 226 -184
rect 234 -191 236 -188
rect 230 -193 236 -191
rect 230 -195 232 -193
rect 234 -195 236 -193
rect 230 -197 236 -195
rect 255 -197 257 -180
rect 269 -184 271 -179
rect 314 -182 316 -177
rect 269 -193 271 -190
rect 269 -195 276 -193
rect 269 -197 272 -195
rect 274 -197 276 -195
rect 223 -203 229 -201
rect 213 -205 219 -203
rect 213 -207 215 -205
rect 217 -207 219 -205
rect 223 -205 225 -203
rect 227 -205 229 -203
rect 223 -207 229 -205
rect 213 -209 219 -207
rect 217 -212 219 -209
rect 224 -212 226 -207
rect 234 -212 236 -197
rect 254 -199 276 -197
rect 254 -202 256 -199
rect 264 -202 266 -199
rect 280 -209 282 -184
rect 287 -187 289 -184
rect 286 -189 292 -187
rect 286 -191 288 -189
rect 290 -191 292 -189
rect 286 -193 292 -191
rect 297 -197 299 -184
rect 276 -211 282 -209
rect 276 -213 278 -211
rect 280 -213 282 -211
rect 254 -219 256 -214
rect 264 -219 266 -214
rect 276 -215 282 -213
rect 280 -218 282 -215
rect 287 -199 299 -197
rect 287 -218 289 -199
rect 304 -201 306 -184
rect 314 -191 316 -188
rect 310 -193 316 -191
rect 310 -195 312 -193
rect 314 -195 316 -193
rect 310 -197 316 -195
rect 303 -203 309 -201
rect 293 -205 299 -203
rect 293 -207 295 -205
rect 297 -207 299 -205
rect 303 -205 305 -203
rect 307 -205 309 -203
rect 303 -207 309 -205
rect 293 -209 299 -207
rect 297 -212 299 -209
rect 304 -212 306 -207
rect 314 -212 316 -197
rect 40 -229 42 -224
rect 47 -232 49 -224
rect 57 -228 59 -224
rect 64 -228 66 -224
rect 74 -232 76 -224
rect 47 -234 76 -232
rect 120 -229 122 -224
rect 127 -232 129 -224
rect 137 -228 139 -224
rect 144 -228 146 -224
rect 154 -232 156 -224
rect 127 -234 156 -232
rect 200 -229 202 -224
rect 207 -232 209 -224
rect 217 -228 219 -224
rect 224 -228 226 -224
rect 234 -232 236 -224
rect 207 -234 236 -232
rect 280 -229 282 -224
rect 287 -232 289 -224
rect 297 -228 299 -224
rect 304 -228 306 -224
rect 314 -232 316 -224
rect 287 -234 316 -232
<< ndif >>
rect -129 27 -122 29
rect -129 25 -127 27
rect -125 25 -122 27
rect -129 23 -122 25
rect -120 27 -113 29
rect -120 25 -117 27
rect -115 25 -113 27
rect -120 23 -113 25
rect -67 24 -60 26
rect -67 22 -65 24
rect -63 22 -60 24
rect -67 20 -60 22
rect -58 23 -50 26
rect -58 20 -48 23
rect -56 14 -48 20
rect -46 14 -41 23
rect -39 21 -32 23
rect -39 19 -36 21
rect -34 19 -32 21
rect -39 17 -32 19
rect 7 21 13 23
rect 22 29 29 31
rect 22 27 24 29
rect 26 27 29 29
rect 22 25 29 27
rect 31 29 38 31
rect 31 27 34 29
rect 36 27 38 29
rect 31 25 38 27
rect 68 25 74 29
rect 7 19 9 21
rect 11 19 15 21
rect 7 17 15 19
rect -39 14 -34 17
rect 10 15 15 17
rect 17 19 24 21
rect 33 19 40 25
rect 42 19 47 25
rect 49 23 57 25
rect 49 21 52 23
rect 54 21 57 23
rect 49 19 57 21
rect 59 19 64 25
rect 66 23 74 25
rect 76 27 83 29
rect 76 25 79 27
rect 81 25 83 27
rect 76 23 83 25
rect 66 19 72 23
rect 17 17 20 19
rect 22 17 24 19
rect 17 15 24 17
rect -56 12 -50 14
rect -56 10 -54 12
rect -52 10 -50 12
rect -56 8 -50 10
rect 68 16 72 19
rect 89 21 95 23
rect 104 29 111 31
rect 104 27 106 29
rect 108 27 111 29
rect 104 25 111 27
rect 113 29 120 31
rect 113 27 116 29
rect 118 27 120 29
rect 113 25 120 27
rect 150 25 156 29
rect 89 19 91 21
rect 93 19 97 21
rect 89 17 97 19
rect 68 12 74 16
rect 92 15 97 17
rect 99 19 106 21
rect 115 19 122 25
rect 124 19 129 25
rect 131 23 139 25
rect 131 21 134 23
rect 136 21 139 23
rect 131 19 139 21
rect 141 19 146 25
rect 148 23 156 25
rect 158 27 165 29
rect 158 25 161 27
rect 163 25 165 27
rect 158 23 165 25
rect 148 19 154 23
rect 99 17 102 19
rect 104 17 106 19
rect 99 15 106 17
rect 68 10 70 12
rect 72 10 74 12
rect 150 16 154 19
rect 170 21 176 23
rect 185 29 192 31
rect 185 27 187 29
rect 189 27 192 29
rect 185 25 192 27
rect 194 29 201 31
rect 194 27 197 29
rect 199 27 201 29
rect 194 25 201 27
rect 231 25 237 29
rect 170 19 172 21
rect 174 19 178 21
rect 170 17 178 19
rect 68 8 74 10
rect 150 12 156 16
rect 173 15 178 17
rect 180 19 187 21
rect 196 19 203 25
rect 205 19 210 25
rect 212 23 220 25
rect 212 21 215 23
rect 217 21 220 23
rect 212 19 220 21
rect 222 19 227 25
rect 229 23 237 25
rect 239 27 246 29
rect 239 25 242 27
rect 244 25 246 27
rect 239 23 246 25
rect 229 19 235 23
rect 180 17 183 19
rect 185 17 187 19
rect 180 15 187 17
rect 150 10 152 12
rect 154 10 156 12
rect 231 16 235 19
rect 253 21 259 23
rect 268 29 275 31
rect 268 27 270 29
rect 272 27 275 29
rect 268 25 275 27
rect 277 29 284 31
rect 277 27 280 29
rect 282 27 284 29
rect 277 25 284 27
rect 314 25 320 29
rect 253 19 255 21
rect 257 19 261 21
rect 253 17 261 19
rect 150 8 156 10
rect 231 12 237 16
rect 256 15 261 17
rect 263 19 270 21
rect 279 19 286 25
rect 288 19 293 25
rect 295 23 303 25
rect 295 21 298 23
rect 300 21 303 23
rect 295 19 303 21
rect 305 19 310 25
rect 312 23 320 25
rect 322 27 329 29
rect 322 25 325 27
rect 327 25 329 27
rect 322 23 329 25
rect 312 19 318 23
rect 263 17 266 19
rect 268 17 270 19
rect 263 15 270 17
rect 231 10 233 12
rect 235 10 237 12
rect 314 16 318 19
rect 231 8 237 10
rect 314 12 320 16
rect 314 10 316 12
rect 318 10 320 12
rect 314 8 320 10
rect -55 -7 -49 -5
rect -55 -9 -53 -7
rect -51 -9 -49 -7
rect -55 -11 -49 -9
rect -55 -17 -47 -11
rect -66 -19 -59 -17
rect -66 -21 -64 -19
rect -62 -21 -59 -19
rect -66 -23 -59 -21
rect -57 -20 -47 -17
rect -45 -20 -40 -11
rect -38 -14 -33 -11
rect 68 -9 74 -7
rect 68 -11 70 -9
rect 72 -11 74 -9
rect -38 -16 -31 -14
rect 10 -16 15 -14
rect -38 -18 -35 -16
rect -33 -18 -31 -16
rect -38 -20 -31 -18
rect 7 -18 15 -16
rect 7 -20 9 -18
rect 11 -20 15 -18
rect 17 -16 24 -14
rect 17 -18 20 -16
rect 22 -18 24 -16
rect 68 -15 74 -11
rect 148 -9 154 -7
rect 148 -11 150 -9
rect 152 -11 154 -9
rect 68 -18 72 -15
rect 90 -16 95 -14
rect 17 -20 24 -18
rect -57 -23 -49 -20
rect -129 -26 -122 -24
rect -129 -28 -127 -26
rect -125 -28 -122 -26
rect -129 -30 -122 -28
rect -120 -26 -113 -24
rect -120 -28 -117 -26
rect -115 -28 -113 -26
rect -120 -30 -113 -28
rect 7 -22 13 -20
rect 33 -24 40 -18
rect 42 -24 47 -18
rect 49 -20 57 -18
rect 49 -22 52 -20
rect 54 -22 57 -20
rect 49 -24 57 -22
rect 59 -24 64 -18
rect 66 -22 72 -18
rect 87 -18 95 -16
rect 87 -20 89 -18
rect 91 -20 95 -18
rect 97 -16 104 -14
rect 97 -18 100 -16
rect 102 -18 104 -16
rect 148 -15 154 -11
rect 231 -9 237 -7
rect 231 -11 233 -9
rect 235 -11 237 -9
rect 148 -18 152 -15
rect 173 -16 178 -14
rect 97 -20 104 -18
rect 87 -22 93 -20
rect 66 -24 74 -22
rect 22 -26 29 -24
rect 22 -28 24 -26
rect 26 -28 29 -26
rect 22 -30 29 -28
rect 31 -26 38 -24
rect 31 -28 34 -26
rect 36 -28 38 -26
rect 31 -30 38 -28
rect 68 -28 74 -24
rect 76 -24 83 -22
rect 76 -26 79 -24
rect 81 -26 83 -24
rect 76 -28 83 -26
rect 113 -24 120 -18
rect 122 -24 127 -18
rect 129 -20 137 -18
rect 129 -22 132 -20
rect 134 -22 137 -20
rect 129 -24 137 -22
rect 139 -24 144 -18
rect 146 -22 152 -18
rect 170 -18 178 -16
rect 170 -20 172 -18
rect 174 -20 178 -18
rect 180 -16 187 -14
rect 180 -18 183 -16
rect 185 -18 187 -16
rect 231 -15 237 -11
rect 311 -9 317 -7
rect 311 -11 313 -9
rect 315 -11 317 -9
rect 231 -18 235 -15
rect 253 -16 258 -14
rect 180 -20 187 -18
rect 170 -22 176 -20
rect 146 -24 154 -22
rect 102 -26 109 -24
rect 102 -28 104 -26
rect 106 -28 109 -26
rect 102 -30 109 -28
rect 111 -26 118 -24
rect 111 -28 114 -26
rect 116 -28 118 -26
rect 111 -30 118 -28
rect 148 -28 154 -24
rect 156 -24 163 -22
rect 156 -26 159 -24
rect 161 -26 163 -24
rect 156 -28 163 -26
rect 196 -24 203 -18
rect 205 -24 210 -18
rect 212 -20 220 -18
rect 212 -22 215 -20
rect 217 -22 220 -20
rect 212 -24 220 -22
rect 222 -24 227 -18
rect 229 -22 235 -18
rect 250 -18 258 -16
rect 250 -20 252 -18
rect 254 -20 258 -18
rect 260 -16 267 -14
rect 260 -18 263 -16
rect 265 -18 267 -16
rect 311 -15 317 -11
rect 311 -18 315 -15
rect 260 -20 267 -18
rect 250 -22 256 -20
rect 229 -24 237 -22
rect 185 -26 192 -24
rect 185 -28 187 -26
rect 189 -28 192 -26
rect 185 -30 192 -28
rect 194 -26 201 -24
rect 194 -28 197 -26
rect 199 -28 201 -26
rect 194 -30 201 -28
rect 231 -28 237 -24
rect 239 -24 246 -22
rect 239 -26 242 -24
rect 244 -26 246 -24
rect 239 -28 246 -26
rect 276 -24 283 -18
rect 285 -24 290 -18
rect 292 -20 300 -18
rect 292 -22 295 -20
rect 297 -22 300 -20
rect 292 -24 300 -22
rect 302 -24 307 -18
rect 309 -22 315 -18
rect 309 -24 317 -22
rect 265 -26 272 -24
rect 265 -28 267 -26
rect 269 -28 272 -26
rect 265 -30 272 -28
rect 274 -26 281 -24
rect 274 -28 277 -26
rect 279 -28 281 -26
rect 274 -30 281 -28
rect 311 -28 317 -24
rect 319 -24 326 -22
rect 319 -26 322 -24
rect 324 -26 326 -24
rect 319 -28 326 -26
rect -65 -134 -58 -132
rect -65 -136 -63 -134
rect -61 -136 -58 -134
rect -65 -138 -58 -136
rect -56 -135 -48 -132
rect -56 -138 -46 -135
rect -54 -144 -46 -138
rect -44 -144 -39 -135
rect -37 -137 -30 -135
rect -37 -139 -34 -137
rect -32 -139 -30 -137
rect -37 -141 -30 -139
rect -37 -144 -32 -141
rect 7 -142 13 -140
rect 22 -134 29 -132
rect 22 -136 24 -134
rect 26 -136 29 -134
rect 22 -138 29 -136
rect 31 -134 38 -132
rect 31 -136 34 -134
rect 36 -136 38 -134
rect 31 -138 38 -136
rect 68 -138 74 -134
rect 7 -144 9 -142
rect 11 -144 15 -142
rect -54 -146 -48 -144
rect -54 -148 -52 -146
rect -50 -148 -48 -146
rect -54 -150 -48 -148
rect 7 -146 15 -144
rect 10 -148 15 -146
rect 17 -144 24 -142
rect 33 -144 40 -138
rect 42 -144 47 -138
rect 49 -140 57 -138
rect 49 -142 52 -140
rect 54 -142 57 -140
rect 49 -144 57 -142
rect 59 -144 64 -138
rect 66 -140 74 -138
rect 76 -136 83 -134
rect 76 -138 79 -136
rect 81 -138 83 -136
rect 76 -140 83 -138
rect 66 -144 72 -140
rect 17 -146 20 -144
rect 22 -146 24 -144
rect 17 -148 24 -146
rect 68 -147 72 -144
rect 87 -142 93 -140
rect 102 -134 109 -132
rect 102 -136 104 -134
rect 106 -136 109 -134
rect 102 -138 109 -136
rect 111 -134 118 -132
rect 111 -136 114 -134
rect 116 -136 118 -134
rect 111 -138 118 -136
rect 148 -138 154 -134
rect 87 -144 89 -142
rect 91 -144 95 -142
rect 87 -146 95 -144
rect 68 -151 74 -147
rect 90 -148 95 -146
rect 97 -144 104 -142
rect 113 -144 120 -138
rect 122 -144 127 -138
rect 129 -140 137 -138
rect 129 -142 132 -140
rect 134 -142 137 -140
rect 129 -144 137 -142
rect 139 -144 144 -138
rect 146 -140 154 -138
rect 156 -136 163 -134
rect 156 -138 159 -136
rect 161 -138 163 -136
rect 156 -140 163 -138
rect 146 -144 152 -140
rect 97 -146 100 -144
rect 102 -146 104 -144
rect 97 -148 104 -146
rect 68 -153 70 -151
rect 72 -153 74 -151
rect 148 -147 152 -144
rect 167 -142 173 -140
rect 182 -134 189 -132
rect 182 -136 184 -134
rect 186 -136 189 -134
rect 182 -138 189 -136
rect 191 -134 198 -132
rect 191 -136 194 -134
rect 196 -136 198 -134
rect 191 -138 198 -136
rect 228 -138 234 -134
rect 167 -144 169 -142
rect 171 -144 175 -142
rect 167 -146 175 -144
rect 68 -155 74 -153
rect 148 -151 154 -147
rect 170 -148 175 -146
rect 177 -144 184 -142
rect 193 -144 200 -138
rect 202 -144 207 -138
rect 209 -140 217 -138
rect 209 -142 212 -140
rect 214 -142 217 -140
rect 209 -144 217 -142
rect 219 -144 224 -138
rect 226 -140 234 -138
rect 236 -136 243 -134
rect 236 -138 239 -136
rect 241 -138 243 -136
rect 236 -140 243 -138
rect 226 -144 232 -140
rect 177 -146 180 -144
rect 182 -146 184 -144
rect 177 -148 184 -146
rect 148 -153 150 -151
rect 152 -153 154 -151
rect 228 -147 232 -144
rect 247 -142 253 -140
rect 262 -134 269 -132
rect 262 -136 264 -134
rect 266 -136 269 -134
rect 262 -138 269 -136
rect 271 -134 278 -132
rect 271 -136 274 -134
rect 276 -136 278 -134
rect 271 -138 278 -136
rect 308 -138 314 -134
rect 247 -144 249 -142
rect 251 -144 255 -142
rect 247 -146 255 -144
rect 148 -155 154 -153
rect 228 -151 234 -147
rect 250 -148 255 -146
rect 257 -144 264 -142
rect 273 -144 280 -138
rect 282 -144 287 -138
rect 289 -140 297 -138
rect 289 -142 292 -140
rect 294 -142 297 -140
rect 289 -144 297 -142
rect 299 -144 304 -138
rect 306 -140 314 -138
rect 316 -136 323 -134
rect 316 -138 319 -136
rect 321 -138 323 -136
rect 316 -140 323 -138
rect 306 -144 312 -140
rect 257 -146 260 -144
rect 262 -146 264 -144
rect 257 -148 264 -146
rect 228 -153 230 -151
rect 232 -153 234 -151
rect 308 -147 312 -144
rect 228 -155 234 -153
rect 308 -151 314 -147
rect 308 -153 310 -151
rect 312 -153 314 -151
rect 308 -155 314 -153
rect -54 -168 -48 -166
rect -54 -170 -52 -168
rect -50 -170 -48 -168
rect -54 -172 -48 -170
rect -54 -178 -46 -172
rect -65 -180 -58 -178
rect -65 -182 -63 -180
rect -61 -182 -58 -180
rect -65 -184 -58 -182
rect -56 -181 -46 -178
rect -44 -181 -39 -172
rect -37 -175 -32 -172
rect 68 -169 74 -167
rect 68 -171 70 -169
rect 72 -171 74 -169
rect -37 -177 -30 -175
rect 10 -176 15 -174
rect -37 -179 -34 -177
rect -32 -179 -30 -177
rect -37 -181 -30 -179
rect 7 -178 15 -176
rect 7 -180 9 -178
rect 11 -180 15 -178
rect 17 -176 24 -174
rect 17 -178 20 -176
rect 22 -178 24 -176
rect 68 -175 74 -171
rect 148 -169 154 -167
rect 148 -171 150 -169
rect 152 -171 154 -169
rect 68 -178 72 -175
rect 90 -176 95 -174
rect 17 -180 24 -178
rect -56 -184 -48 -181
rect 7 -182 13 -180
rect 33 -184 40 -178
rect 42 -184 47 -178
rect 49 -180 57 -178
rect 49 -182 52 -180
rect 54 -182 57 -180
rect 49 -184 57 -182
rect 59 -184 64 -178
rect 66 -182 72 -178
rect 87 -178 95 -176
rect 87 -180 89 -178
rect 91 -180 95 -178
rect 97 -176 104 -174
rect 97 -178 100 -176
rect 102 -178 104 -176
rect 148 -175 154 -171
rect 228 -169 234 -167
rect 228 -171 230 -169
rect 232 -171 234 -169
rect 148 -178 152 -175
rect 170 -176 175 -174
rect 97 -180 104 -178
rect 87 -182 93 -180
rect 66 -184 74 -182
rect 22 -186 29 -184
rect 22 -188 24 -186
rect 26 -188 29 -186
rect 22 -190 29 -188
rect 31 -186 38 -184
rect 31 -188 34 -186
rect 36 -188 38 -186
rect 31 -190 38 -188
rect 68 -188 74 -184
rect 76 -184 83 -182
rect 76 -186 79 -184
rect 81 -186 83 -184
rect 76 -188 83 -186
rect 113 -184 120 -178
rect 122 -184 127 -178
rect 129 -180 137 -178
rect 129 -182 132 -180
rect 134 -182 137 -180
rect 129 -184 137 -182
rect 139 -184 144 -178
rect 146 -182 152 -178
rect 167 -178 175 -176
rect 167 -180 169 -178
rect 171 -180 175 -178
rect 177 -176 184 -174
rect 177 -178 180 -176
rect 182 -178 184 -176
rect 228 -175 234 -171
rect 308 -169 314 -167
rect 308 -171 310 -169
rect 312 -171 314 -169
rect 228 -178 232 -175
rect 250 -176 255 -174
rect 177 -180 184 -178
rect 167 -182 173 -180
rect 146 -184 154 -182
rect 102 -186 109 -184
rect 102 -188 104 -186
rect 106 -188 109 -186
rect 102 -190 109 -188
rect 111 -186 118 -184
rect 111 -188 114 -186
rect 116 -188 118 -186
rect 111 -190 118 -188
rect 148 -188 154 -184
rect 156 -184 163 -182
rect 156 -186 159 -184
rect 161 -186 163 -184
rect 156 -188 163 -186
rect 193 -184 200 -178
rect 202 -184 207 -178
rect 209 -180 217 -178
rect 209 -182 212 -180
rect 214 -182 217 -180
rect 209 -184 217 -182
rect 219 -184 224 -178
rect 226 -182 232 -178
rect 247 -178 255 -176
rect 247 -180 249 -178
rect 251 -180 255 -178
rect 257 -176 264 -174
rect 257 -178 260 -176
rect 262 -178 264 -176
rect 308 -175 314 -171
rect 308 -178 312 -175
rect 257 -180 264 -178
rect 247 -182 253 -180
rect 226 -184 234 -182
rect 182 -186 189 -184
rect 182 -188 184 -186
rect 186 -188 189 -186
rect 182 -190 189 -188
rect 191 -186 198 -184
rect 191 -188 194 -186
rect 196 -188 198 -186
rect 191 -190 198 -188
rect 228 -188 234 -184
rect 236 -184 243 -182
rect 236 -186 239 -184
rect 241 -186 243 -184
rect 236 -188 243 -186
rect 273 -184 280 -178
rect 282 -184 287 -178
rect 289 -180 297 -178
rect 289 -182 292 -180
rect 294 -182 297 -180
rect 289 -184 297 -182
rect 299 -184 304 -178
rect 306 -182 312 -178
rect 306 -184 314 -182
rect 262 -186 269 -184
rect 262 -188 264 -186
rect 266 -188 269 -186
rect 262 -190 269 -188
rect 271 -186 278 -184
rect 271 -188 274 -186
rect 276 -188 278 -186
rect 271 -190 278 -188
rect 308 -188 314 -184
rect 316 -184 323 -182
rect 316 -186 319 -184
rect 321 -186 323 -184
rect 316 -188 323 -186
<< pdif >>
rect -129 70 -123 72
rect -129 68 -127 70
rect -125 68 -123 70
rect -129 64 -123 68
rect -129 53 -124 64
rect 33 63 40 65
rect 33 61 35 63
rect 37 61 40 63
rect -129 41 -122 53
rect -120 47 -115 53
rect -65 49 -60 55
rect -67 47 -60 49
rect -120 45 -113 47
rect -120 43 -117 45
rect -115 43 -113 45
rect -67 45 -65 47
rect -63 45 -60 47
rect -67 43 -60 45
rect -58 53 -52 55
rect 33 59 40 61
rect 42 59 47 65
rect 49 63 57 65
rect 49 61 52 63
rect 54 61 57 63
rect 49 59 57 61
rect -58 47 -50 53
rect -58 45 -55 47
rect -53 45 -50 47
rect -58 43 -50 45
rect -48 47 -40 53
rect -48 45 -45 47
rect -43 45 -40 47
rect -48 43 -40 45
rect -38 51 -31 53
rect -38 49 -35 51
rect -33 49 -31 51
rect 9 49 14 55
rect -38 43 -31 49
rect 7 47 14 49
rect 7 45 9 47
rect 11 45 14 47
rect 7 43 14 45
rect 16 53 24 55
rect 16 51 19 53
rect 21 51 24 53
rect 16 43 24 51
rect 26 53 33 55
rect 26 51 29 53
rect 31 51 33 53
rect 26 49 33 51
rect 26 43 31 49
rect -120 41 -113 43
rect 52 53 57 59
rect 59 53 64 65
rect 66 63 74 65
rect 66 61 69 63
rect 71 61 74 63
rect 66 53 74 61
rect 76 59 81 65
rect 115 63 122 65
rect 115 61 117 63
rect 119 61 122 63
rect 76 57 83 59
rect 76 55 79 57
rect 81 55 83 57
rect 115 59 122 61
rect 124 59 129 65
rect 131 63 139 65
rect 131 61 134 63
rect 136 61 139 63
rect 131 59 139 61
rect 76 53 83 55
rect 91 49 96 55
rect 89 47 96 49
rect 89 45 91 47
rect 93 45 96 47
rect 89 43 96 45
rect 98 53 106 55
rect 98 51 101 53
rect 103 51 106 53
rect 98 43 106 51
rect 108 53 115 55
rect 108 51 111 53
rect 113 51 115 53
rect 108 49 115 51
rect 108 43 113 49
rect 134 53 139 59
rect 141 53 146 65
rect 148 63 156 65
rect 148 61 151 63
rect 153 61 156 63
rect 148 53 156 61
rect 158 59 163 65
rect 196 63 203 65
rect 196 61 198 63
rect 200 61 203 63
rect 158 57 165 59
rect 158 55 161 57
rect 163 55 165 57
rect 196 59 203 61
rect 205 59 210 65
rect 212 63 220 65
rect 212 61 215 63
rect 217 61 220 63
rect 212 59 220 61
rect 158 53 165 55
rect 172 49 177 55
rect 170 47 177 49
rect 170 45 172 47
rect 174 45 177 47
rect 170 43 177 45
rect 179 53 187 55
rect 179 51 182 53
rect 184 51 187 53
rect 179 43 187 51
rect 189 53 196 55
rect 189 51 192 53
rect 194 51 196 53
rect 189 49 196 51
rect 189 43 194 49
rect 215 53 220 59
rect 222 53 227 65
rect 229 63 237 65
rect 229 61 232 63
rect 234 61 237 63
rect 229 53 237 61
rect 239 59 244 65
rect 279 63 286 65
rect 279 61 281 63
rect 283 61 286 63
rect 239 57 246 59
rect 239 55 242 57
rect 244 55 246 57
rect 279 59 286 61
rect 288 59 293 65
rect 295 63 303 65
rect 295 61 298 63
rect 300 61 303 63
rect 295 59 303 61
rect 239 53 246 55
rect 255 49 260 55
rect 253 47 260 49
rect 253 45 255 47
rect 257 45 260 47
rect 253 43 260 45
rect 262 53 270 55
rect 262 51 265 53
rect 267 51 270 53
rect 262 43 270 51
rect 272 53 279 55
rect 272 51 275 53
rect 277 51 279 53
rect 272 49 279 51
rect 272 43 277 49
rect 298 53 303 59
rect 305 53 310 65
rect 312 63 320 65
rect 312 61 315 63
rect 317 61 320 63
rect 312 53 320 61
rect 322 59 327 65
rect 322 57 329 59
rect 322 55 325 57
rect 327 55 329 57
rect 322 53 329 55
rect -66 -42 -59 -40
rect -129 -54 -122 -42
rect -120 -44 -113 -42
rect -120 -46 -117 -44
rect -115 -46 -113 -44
rect -66 -44 -64 -42
rect -62 -44 -59 -42
rect -66 -46 -59 -44
rect -120 -48 -113 -46
rect -120 -54 -115 -48
rect -64 -52 -59 -46
rect -57 -42 -49 -40
rect -57 -44 -54 -42
rect -52 -44 -49 -42
rect -57 -50 -49 -44
rect -47 -42 -39 -40
rect -47 -44 -44 -42
rect -42 -44 -39 -42
rect -47 -50 -39 -44
rect -37 -46 -30 -40
rect -37 -48 -34 -46
rect -32 -48 -30 -46
rect 7 -44 14 -42
rect 7 -46 9 -44
rect 11 -46 14 -44
rect 7 -48 14 -46
rect -37 -50 -30 -48
rect -57 -52 -51 -50
rect -129 -65 -124 -54
rect 9 -54 14 -48
rect 16 -50 24 -42
rect 16 -52 19 -50
rect 21 -52 24 -50
rect 16 -54 24 -52
rect 26 -48 31 -42
rect 26 -50 33 -48
rect 26 -52 29 -50
rect 31 -52 33 -50
rect 26 -54 33 -52
rect 87 -44 94 -42
rect 87 -46 89 -44
rect 91 -46 94 -44
rect 87 -48 94 -46
rect 52 -58 57 -52
rect 33 -60 40 -58
rect 33 -62 35 -60
rect 37 -62 40 -60
rect 33 -64 40 -62
rect 42 -64 47 -58
rect 49 -60 57 -58
rect 49 -62 52 -60
rect 54 -62 57 -60
rect 49 -64 57 -62
rect 59 -64 64 -52
rect 66 -60 74 -52
rect 66 -62 69 -60
rect 71 -62 74 -60
rect 66 -64 74 -62
rect 76 -54 83 -52
rect 89 -54 94 -48
rect 96 -50 104 -42
rect 96 -52 99 -50
rect 101 -52 104 -50
rect 96 -54 104 -52
rect 106 -48 111 -42
rect 106 -50 113 -48
rect 106 -52 109 -50
rect 111 -52 113 -50
rect 106 -54 113 -52
rect 76 -56 79 -54
rect 81 -56 83 -54
rect 76 -58 83 -56
rect 76 -64 81 -58
rect 170 -44 177 -42
rect 170 -46 172 -44
rect 174 -46 177 -44
rect 170 -48 177 -46
rect 132 -58 137 -52
rect 113 -60 120 -58
rect 113 -62 115 -60
rect 117 -62 120 -60
rect 113 -64 120 -62
rect 122 -64 127 -58
rect 129 -60 137 -58
rect 129 -62 132 -60
rect 134 -62 137 -60
rect 129 -64 137 -62
rect 139 -64 144 -52
rect 146 -60 154 -52
rect 146 -62 149 -60
rect 151 -62 154 -60
rect 146 -64 154 -62
rect 156 -54 163 -52
rect 172 -54 177 -48
rect 179 -50 187 -42
rect 179 -52 182 -50
rect 184 -52 187 -50
rect 179 -54 187 -52
rect 189 -48 194 -42
rect 189 -50 196 -48
rect 189 -52 192 -50
rect 194 -52 196 -50
rect 189 -54 196 -52
rect 156 -56 159 -54
rect 161 -56 163 -54
rect 156 -58 163 -56
rect 156 -64 161 -58
rect 250 -44 257 -42
rect 250 -46 252 -44
rect 254 -46 257 -44
rect 250 -48 257 -46
rect 215 -58 220 -52
rect 196 -60 203 -58
rect 196 -62 198 -60
rect 200 -62 203 -60
rect 196 -64 203 -62
rect 205 -64 210 -58
rect 212 -60 220 -58
rect 212 -62 215 -60
rect 217 -62 220 -60
rect 212 -64 220 -62
rect 222 -64 227 -52
rect 229 -60 237 -52
rect 229 -62 232 -60
rect 234 -62 237 -60
rect 229 -64 237 -62
rect 239 -54 246 -52
rect 252 -54 257 -48
rect 259 -50 267 -42
rect 259 -52 262 -50
rect 264 -52 267 -50
rect 259 -54 267 -52
rect 269 -48 274 -42
rect 269 -50 276 -48
rect 269 -52 272 -50
rect 274 -52 276 -50
rect 269 -54 276 -52
rect 239 -56 242 -54
rect 244 -56 246 -54
rect 239 -58 246 -56
rect 239 -64 244 -58
rect 295 -58 300 -52
rect 276 -60 283 -58
rect 276 -62 278 -60
rect 280 -62 283 -60
rect 276 -64 283 -62
rect 285 -64 290 -58
rect 292 -60 300 -58
rect 292 -62 295 -60
rect 297 -62 300 -60
rect 292 -64 300 -62
rect 302 -64 307 -52
rect 309 -60 317 -52
rect 309 -62 312 -60
rect 314 -62 317 -60
rect 309 -64 317 -62
rect 319 -54 326 -52
rect 319 -56 322 -54
rect 324 -56 326 -54
rect 319 -58 326 -56
rect 319 -64 324 -58
rect -129 -69 -123 -65
rect -129 -71 -127 -69
rect -125 -71 -123 -69
rect -129 -73 -123 -71
rect 33 -100 40 -98
rect -63 -109 -58 -103
rect -65 -111 -58 -109
rect -65 -113 -63 -111
rect -61 -113 -58 -111
rect -65 -115 -58 -113
rect -56 -105 -50 -103
rect 33 -102 35 -100
rect 37 -102 40 -100
rect -56 -111 -48 -105
rect -56 -113 -53 -111
rect -51 -113 -48 -111
rect -56 -115 -48 -113
rect -46 -111 -38 -105
rect -46 -113 -43 -111
rect -41 -113 -38 -111
rect -46 -115 -38 -113
rect -36 -107 -29 -105
rect -36 -109 -33 -107
rect -31 -109 -29 -107
rect 33 -104 40 -102
rect 42 -104 47 -98
rect 49 -100 57 -98
rect 49 -102 52 -100
rect 54 -102 57 -100
rect 49 -104 57 -102
rect -36 -115 -29 -109
rect 9 -114 14 -108
rect 7 -116 14 -114
rect 7 -118 9 -116
rect 11 -118 14 -116
rect 7 -120 14 -118
rect 16 -110 24 -108
rect 16 -112 19 -110
rect 21 -112 24 -110
rect 16 -120 24 -112
rect 26 -110 33 -108
rect 26 -112 29 -110
rect 31 -112 33 -110
rect 26 -114 33 -112
rect 26 -120 31 -114
rect 52 -110 57 -104
rect 59 -110 64 -98
rect 66 -100 74 -98
rect 66 -102 69 -100
rect 71 -102 74 -100
rect 66 -110 74 -102
rect 76 -104 81 -98
rect 113 -100 120 -98
rect 113 -102 115 -100
rect 117 -102 120 -100
rect 76 -106 83 -104
rect 76 -108 79 -106
rect 81 -108 83 -106
rect 113 -104 120 -102
rect 122 -104 127 -98
rect 129 -100 137 -98
rect 129 -102 132 -100
rect 134 -102 137 -100
rect 129 -104 137 -102
rect 76 -110 83 -108
rect 89 -114 94 -108
rect 87 -116 94 -114
rect 87 -118 89 -116
rect 91 -118 94 -116
rect 87 -120 94 -118
rect 96 -110 104 -108
rect 96 -112 99 -110
rect 101 -112 104 -110
rect 96 -120 104 -112
rect 106 -110 113 -108
rect 106 -112 109 -110
rect 111 -112 113 -110
rect 106 -114 113 -112
rect 106 -120 111 -114
rect 132 -110 137 -104
rect 139 -110 144 -98
rect 146 -100 154 -98
rect 146 -102 149 -100
rect 151 -102 154 -100
rect 146 -110 154 -102
rect 156 -104 161 -98
rect 193 -100 200 -98
rect 193 -102 195 -100
rect 197 -102 200 -100
rect 156 -106 163 -104
rect 156 -108 159 -106
rect 161 -108 163 -106
rect 193 -104 200 -102
rect 202 -104 207 -98
rect 209 -100 217 -98
rect 209 -102 212 -100
rect 214 -102 217 -100
rect 209 -104 217 -102
rect 156 -110 163 -108
rect 169 -114 174 -108
rect 167 -116 174 -114
rect 167 -118 169 -116
rect 171 -118 174 -116
rect 167 -120 174 -118
rect 176 -110 184 -108
rect 176 -112 179 -110
rect 181 -112 184 -110
rect 176 -120 184 -112
rect 186 -110 193 -108
rect 186 -112 189 -110
rect 191 -112 193 -110
rect 186 -114 193 -112
rect 186 -120 191 -114
rect 212 -110 217 -104
rect 219 -110 224 -98
rect 226 -100 234 -98
rect 226 -102 229 -100
rect 231 -102 234 -100
rect 226 -110 234 -102
rect 236 -104 241 -98
rect 273 -100 280 -98
rect 273 -102 275 -100
rect 277 -102 280 -100
rect 236 -106 243 -104
rect 236 -108 239 -106
rect 241 -108 243 -106
rect 273 -104 280 -102
rect 282 -104 287 -98
rect 289 -100 297 -98
rect 289 -102 292 -100
rect 294 -102 297 -100
rect 289 -104 297 -102
rect 236 -110 243 -108
rect 249 -114 254 -108
rect 247 -116 254 -114
rect 247 -118 249 -116
rect 251 -118 254 -116
rect 247 -120 254 -118
rect 256 -110 264 -108
rect 256 -112 259 -110
rect 261 -112 264 -110
rect 256 -120 264 -112
rect 266 -110 273 -108
rect 266 -112 269 -110
rect 271 -112 273 -110
rect 266 -114 273 -112
rect 266 -120 271 -114
rect 292 -110 297 -104
rect 299 -110 304 -98
rect 306 -100 314 -98
rect 306 -102 309 -100
rect 311 -102 314 -100
rect 306 -110 314 -102
rect 316 -104 321 -98
rect 316 -106 323 -104
rect 316 -108 319 -106
rect 321 -108 323 -106
rect 316 -110 323 -108
rect -65 -203 -58 -201
rect -65 -205 -63 -203
rect -61 -205 -58 -203
rect -65 -207 -58 -205
rect -63 -213 -58 -207
rect -56 -203 -48 -201
rect -56 -205 -53 -203
rect -51 -205 -48 -203
rect -56 -211 -48 -205
rect -46 -203 -38 -201
rect -46 -205 -43 -203
rect -41 -205 -38 -203
rect -46 -211 -38 -205
rect -36 -207 -29 -201
rect -36 -209 -33 -207
rect -31 -209 -29 -207
rect 7 -204 14 -202
rect 7 -206 9 -204
rect 11 -206 14 -204
rect 7 -208 14 -206
rect -36 -211 -29 -209
rect -56 -213 -50 -211
rect 9 -214 14 -208
rect 16 -210 24 -202
rect 16 -212 19 -210
rect 21 -212 24 -210
rect 16 -214 24 -212
rect 26 -208 31 -202
rect 26 -210 33 -208
rect 26 -212 29 -210
rect 31 -212 33 -210
rect 26 -214 33 -212
rect 87 -204 94 -202
rect 87 -206 89 -204
rect 91 -206 94 -204
rect 87 -208 94 -206
rect 52 -218 57 -212
rect 33 -220 40 -218
rect 33 -222 35 -220
rect 37 -222 40 -220
rect 33 -224 40 -222
rect 42 -224 47 -218
rect 49 -220 57 -218
rect 49 -222 52 -220
rect 54 -222 57 -220
rect 49 -224 57 -222
rect 59 -224 64 -212
rect 66 -220 74 -212
rect 66 -222 69 -220
rect 71 -222 74 -220
rect 66 -224 74 -222
rect 76 -214 83 -212
rect 89 -214 94 -208
rect 96 -210 104 -202
rect 96 -212 99 -210
rect 101 -212 104 -210
rect 96 -214 104 -212
rect 106 -208 111 -202
rect 106 -210 113 -208
rect 106 -212 109 -210
rect 111 -212 113 -210
rect 106 -214 113 -212
rect 76 -216 79 -214
rect 81 -216 83 -214
rect 76 -218 83 -216
rect 76 -224 81 -218
rect 167 -204 174 -202
rect 167 -206 169 -204
rect 171 -206 174 -204
rect 167 -208 174 -206
rect 132 -218 137 -212
rect 113 -220 120 -218
rect 113 -222 115 -220
rect 117 -222 120 -220
rect 113 -224 120 -222
rect 122 -224 127 -218
rect 129 -220 137 -218
rect 129 -222 132 -220
rect 134 -222 137 -220
rect 129 -224 137 -222
rect 139 -224 144 -212
rect 146 -220 154 -212
rect 146 -222 149 -220
rect 151 -222 154 -220
rect 146 -224 154 -222
rect 156 -214 163 -212
rect 169 -214 174 -208
rect 176 -210 184 -202
rect 176 -212 179 -210
rect 181 -212 184 -210
rect 176 -214 184 -212
rect 186 -208 191 -202
rect 186 -210 193 -208
rect 186 -212 189 -210
rect 191 -212 193 -210
rect 186 -214 193 -212
rect 156 -216 159 -214
rect 161 -216 163 -214
rect 156 -218 163 -216
rect 156 -224 161 -218
rect 247 -204 254 -202
rect 247 -206 249 -204
rect 251 -206 254 -204
rect 247 -208 254 -206
rect 212 -218 217 -212
rect 193 -220 200 -218
rect 193 -222 195 -220
rect 197 -222 200 -220
rect 193 -224 200 -222
rect 202 -224 207 -218
rect 209 -220 217 -218
rect 209 -222 212 -220
rect 214 -222 217 -220
rect 209 -224 217 -222
rect 219 -224 224 -212
rect 226 -220 234 -212
rect 226 -222 229 -220
rect 231 -222 234 -220
rect 226 -224 234 -222
rect 236 -214 243 -212
rect 249 -214 254 -208
rect 256 -210 264 -202
rect 256 -212 259 -210
rect 261 -212 264 -210
rect 256 -214 264 -212
rect 266 -208 271 -202
rect 266 -210 273 -208
rect 266 -212 269 -210
rect 271 -212 273 -210
rect 266 -214 273 -212
rect 236 -216 239 -214
rect 241 -216 243 -214
rect 236 -218 243 -216
rect 236 -224 241 -218
rect 292 -218 297 -212
rect 273 -220 280 -218
rect 273 -222 275 -220
rect 277 -222 280 -220
rect 273 -224 280 -222
rect 282 -224 287 -218
rect 289 -220 297 -218
rect 289 -222 292 -220
rect 294 -222 297 -220
rect 289 -224 297 -222
rect 299 -224 304 -212
rect 306 -220 314 -212
rect 306 -222 309 -220
rect 311 -222 314 -220
rect 306 -224 314 -222
rect 316 -214 323 -212
rect 316 -216 319 -214
rect 321 -216 323 -214
rect 316 -218 323 -216
rect 316 -224 321 -218
<< alu1 >>
rect -71 75 -27 77
rect 3 75 333 77
rect -133 72 333 75
rect -133 71 -64 72
rect -133 70 -105 71
rect -133 68 -127 70
rect -125 68 -117 70
rect -115 68 -105 70
rect -71 70 -64 71
rect -62 70 -50 72
rect -48 70 -36 72
rect -34 71 10 72
rect -34 70 -27 71
rect -71 69 -27 70
rect -133 67 -105 68
rect -97 62 -59 64
rect -55 62 -39 64
rect -150 60 -117 62
rect -150 58 -120 60
rect -118 58 -117 60
rect -150 56 -117 58
rect -97 60 -48 62
rect -46 60 -39 62
rect -150 -17 -146 56
rect -129 48 -125 56
rect -121 45 -113 46
rect -121 43 -117 45
rect -115 43 -113 45
rect -121 42 -113 43
rect -121 38 -117 42
rect -97 41 -93 60
rect -98 38 -93 41
rect -129 37 -93 38
rect -67 47 -63 56
rect -67 45 -65 47
rect -67 38 -63 45
rect -52 58 -39 60
rect -52 51 -46 58
rect -129 35 -101 37
rect -99 35 -94 37
rect -129 34 -94 35
rect -67 36 -66 38
rect -64 36 -63 38
rect -129 32 -117 34
rect -129 27 -123 32
rect -81 29 -77 31
rect -129 25 -127 27
rect -125 25 -123 27
rect -129 24 -123 25
rect -81 27 -80 29
rect -78 27 -77 29
rect -133 10 -105 11
rect -133 8 -126 10
rect -124 8 -118 10
rect -116 9 -88 10
rect -116 8 -91 9
rect -133 7 -91 8
rect -89 7 -88 9
rect -133 6 -88 7
rect -133 3 -105 6
rect -112 -4 -108 3
rect -133 -9 -105 -4
rect -133 -11 -126 -9
rect -124 -11 -118 -9
rect -116 -11 -105 -9
rect -133 -12 -105 -11
rect -164 -18 -89 -17
rect -164 -20 -92 -18
rect -90 -20 -89 -18
rect -164 -21 -89 -20
rect -164 -219 -160 -21
rect -129 -26 -123 -25
rect -129 -28 -127 -26
rect -125 -28 -123 -26
rect -129 -33 -123 -28
rect -81 -25 -77 27
rect -67 24 -63 36
rect -67 22 -65 24
rect -63 22 -55 24
rect -67 18 -55 22
rect -44 31 -40 32
rect -35 31 -31 40
rect -44 30 -31 31
rect -44 28 -39 30
rect -37 28 -31 30
rect -44 26 -31 28
rect -71 12 -26 13
rect -71 10 -64 12
rect -62 10 -54 12
rect -52 10 -26 12
rect -71 8 -29 10
rect -27 8 -26 10
rect -71 5 -26 8
rect -34 -2 -30 5
rect -71 -3 -26 -2
rect -71 -5 -70 -3
rect -68 -5 -26 -3
rect -71 -6 -26 -5
rect -70 -7 -26 -6
rect -70 -9 -63 -7
rect -61 -9 -53 -7
rect -51 -9 -26 -7
rect -70 -10 -26 -9
rect -81 -27 -80 -25
rect -78 -27 -77 -25
rect -81 -30 -77 -27
rect -129 -34 -117 -33
rect -82 -34 -77 -30
rect -66 -19 -54 -15
rect -66 -21 -64 -19
rect -62 -21 -54 -19
rect -66 -34 -62 -21
rect -43 -25 -30 -23
rect -43 -27 -38 -25
rect -36 -27 -30 -25
rect -43 -28 -30 -27
rect -129 -38 -78 -34
rect -66 -36 -65 -34
rect -63 -36 -62 -34
rect -129 -39 -117 -38
rect -121 -43 -117 -39
rect -66 -42 -62 -36
rect -121 -44 -113 -43
rect -121 -46 -117 -44
rect -115 -46 -113 -44
rect -121 -47 -113 -46
rect -66 -44 -64 -42
rect -129 -57 -125 -49
rect -66 -53 -62 -44
rect -34 -37 -30 -28
rect -152 -59 -117 -57
rect -152 -61 -120 -59
rect -118 -61 -117 -59
rect -152 -63 -117 -61
rect -152 -129 -147 -63
rect -51 -55 -45 -48
rect -51 -57 -38 -55
rect -51 -59 -47 -57
rect -45 -59 -38 -57
rect -51 -61 -38 -59
rect -70 -67 -26 -66
rect -133 -69 -105 -68
rect -70 -69 -63 -67
rect -61 -69 -49 -67
rect -47 -69 -35 -67
rect -33 -68 -26 -67
rect -13 -68 -9 71
rect 3 70 10 71
rect 12 70 18 72
rect 20 70 92 72
rect 94 70 100 72
rect 102 70 173 72
rect 175 70 181 72
rect 183 70 256 72
rect 258 70 264 72
rect 266 70 333 72
rect 3 69 333 70
rect 7 47 12 49
rect 7 45 9 47
rect 11 45 12 47
rect 7 43 12 45
rect 7 32 11 43
rect 7 26 19 32
rect 7 21 13 26
rect 7 19 9 21
rect 11 19 13 21
rect 7 18 13 19
rect 63 46 68 48
rect 63 44 65 46
rect 67 44 68 46
rect 63 42 68 44
rect 63 31 67 42
rect 54 27 67 31
rect 71 36 75 38
rect 71 34 72 36
rect 74 34 75 36
rect 71 23 75 34
rect 89 47 94 49
rect 89 45 91 47
rect 93 45 94 47
rect 89 43 94 45
rect 89 32 93 43
rect 89 26 101 32
rect 62 19 75 23
rect 89 21 95 26
rect 89 19 91 21
rect 93 19 95 21
rect 89 18 95 19
rect 145 46 150 48
rect 145 44 147 46
rect 149 44 150 46
rect 145 42 150 44
rect 145 31 149 42
rect 136 27 149 31
rect 153 36 157 38
rect 153 34 154 36
rect 156 34 157 36
rect 153 23 157 34
rect 170 47 175 49
rect 170 45 172 47
rect 174 45 175 47
rect 170 43 175 45
rect 170 32 174 43
rect 170 26 182 32
rect 144 19 157 23
rect 170 21 176 26
rect 170 19 172 21
rect 174 19 176 21
rect 170 18 176 19
rect 226 46 231 48
rect 226 44 228 46
rect 230 44 231 46
rect 226 42 231 44
rect 226 31 230 42
rect 217 27 230 31
rect 234 36 238 38
rect 234 34 235 36
rect 237 34 238 36
rect 234 23 238 34
rect 253 47 258 49
rect 253 45 255 47
rect 257 45 258 47
rect 253 43 258 45
rect 253 32 257 43
rect 253 26 265 32
rect 225 19 238 23
rect 253 21 259 26
rect 253 19 255 21
rect 257 19 259 21
rect 253 18 259 19
rect 309 46 314 48
rect 309 44 311 46
rect 313 44 314 46
rect 309 42 314 44
rect 309 31 313 42
rect 300 27 313 31
rect 317 36 321 38
rect 317 34 318 36
rect 320 34 321 36
rect 317 23 321 34
rect 308 19 321 23
rect 3 12 333 13
rect 3 10 30 12
rect 32 10 70 12
rect 72 10 112 12
rect 114 10 152 12
rect 154 10 193 12
rect 195 10 233 12
rect 235 10 276 12
rect 278 10 316 12
rect 318 10 346 12
rect 3 8 4 10
rect 6 8 346 10
rect 3 5 333 8
rect 56 -4 61 5
rect 3 -9 330 -4
rect 3 -11 30 -9
rect 32 -11 70 -9
rect 72 -11 110 -9
rect 112 -11 150 -9
rect 152 -11 193 -9
rect 195 -11 233 -9
rect 235 -11 273 -9
rect 275 -11 313 -9
rect 315 -11 330 -9
rect 3 -12 330 -11
rect 7 -18 13 -17
rect 7 -20 9 -18
rect 11 -20 13 -18
rect 7 -25 13 -20
rect 7 -31 19 -25
rect 7 -42 11 -31
rect 87 -18 93 -17
rect 62 -22 75 -18
rect 87 -20 89 -18
rect 91 -20 93 -18
rect 54 -30 67 -26
rect 7 -44 12 -42
rect 7 -46 9 -44
rect 11 -46 12 -44
rect 7 -48 12 -46
rect 63 -41 67 -30
rect 71 -33 75 -22
rect 71 -35 72 -33
rect 74 -35 75 -33
rect 71 -37 75 -35
rect 63 -43 68 -41
rect 63 -45 65 -43
rect 67 -45 68 -43
rect 63 -47 68 -45
rect 87 -25 93 -20
rect 87 -31 99 -25
rect 87 -42 91 -31
rect 170 -18 176 -17
rect 142 -22 155 -18
rect 170 -20 172 -18
rect 174 -20 176 -18
rect 134 -30 147 -26
rect 87 -44 92 -42
rect 87 -46 89 -44
rect 91 -46 92 -44
rect 87 -48 92 -46
rect 143 -41 147 -30
rect 151 -33 155 -22
rect 151 -35 152 -33
rect 154 -35 155 -33
rect 151 -37 155 -35
rect 143 -43 148 -41
rect 143 -45 145 -43
rect 147 -45 148 -43
rect 143 -47 148 -45
rect 170 -25 176 -20
rect 170 -31 182 -25
rect 170 -42 174 -31
rect 250 -18 256 -17
rect 225 -22 238 -18
rect 250 -20 252 -18
rect 254 -20 256 -18
rect 217 -30 230 -26
rect 170 -44 175 -42
rect 170 -46 172 -44
rect 174 -46 175 -44
rect 170 -48 175 -46
rect 226 -41 230 -30
rect 234 -33 238 -22
rect 234 -35 235 -33
rect 237 -35 238 -33
rect 234 -37 238 -35
rect 226 -43 231 -41
rect 226 -45 228 -43
rect 230 -45 231 -43
rect 226 -47 231 -45
rect 250 -25 256 -20
rect 250 -31 262 -25
rect 250 -42 254 -31
rect 305 -22 318 -18
rect 297 -30 310 -26
rect 250 -44 255 -42
rect 250 -46 252 -44
rect 254 -46 255 -44
rect 250 -48 255 -46
rect 306 -41 310 -30
rect 314 -33 318 -22
rect 314 -35 315 -33
rect 317 -35 318 -33
rect 314 -37 318 -35
rect 306 -43 311 -41
rect 306 -45 308 -43
rect 310 -45 311 -43
rect 306 -47 311 -45
rect -33 -69 -9 -68
rect -133 -71 -127 -69
rect -125 -71 -117 -69
rect -115 -71 -9 -69
rect -133 -72 -9 -71
rect -133 -73 -26 -72
rect -133 -76 -105 -73
rect -70 -74 -26 -73
rect -64 -81 -60 -74
rect -69 -86 -25 -81
rect -69 -88 -62 -86
rect -60 -88 -48 -86
rect -46 -88 -34 -86
rect -32 -88 -25 -86
rect -69 -89 -25 -88
rect -13 -88 -9 -72
rect 3 -69 330 -68
rect 3 -71 10 -69
rect 12 -71 18 -69
rect 20 -71 90 -69
rect 92 -71 98 -69
rect 100 -71 173 -69
rect 175 -71 181 -69
rect 183 -71 253 -69
rect 255 -71 261 -69
rect 263 -71 330 -69
rect 3 -76 330 -71
rect 162 -86 167 -76
rect 3 -88 327 -86
rect -152 -131 -151 -129
rect -149 -131 -147 -129
rect -152 -186 -147 -131
rect -65 -111 -61 -102
rect -65 -113 -63 -111
rect -65 -119 -61 -113
rect -50 -96 -37 -94
rect -50 -98 -46 -96
rect -44 -98 -37 -96
rect -50 -100 -37 -98
rect -50 -107 -44 -100
rect -13 -91 327 -88
rect -13 -92 10 -91
rect -65 -121 -64 -119
rect -62 -121 -61 -119
rect -65 -134 -61 -121
rect -65 -136 -63 -134
rect -61 -136 -53 -134
rect -65 -140 -53 -136
rect -33 -127 -29 -118
rect -42 -128 -29 -127
rect -42 -130 -37 -128
rect -35 -130 -29 -128
rect -42 -132 -29 -130
rect -69 -146 -25 -145
rect -69 -148 -62 -146
rect -60 -148 -52 -146
rect -50 -148 -25 -146
rect -69 -153 -25 -148
rect -37 -163 -33 -153
rect -69 -165 -24 -163
rect -69 -167 -27 -165
rect -25 -167 -24 -165
rect -69 -168 -24 -167
rect -69 -170 -62 -168
rect -60 -170 -52 -168
rect -50 -170 -24 -168
rect -69 -171 -24 -170
rect -152 -188 -151 -186
rect -149 -188 -147 -186
rect -152 -189 -147 -188
rect -65 -180 -53 -176
rect -65 -182 -63 -180
rect -61 -182 -53 -180
rect -65 -203 -61 -182
rect -42 -186 -29 -184
rect -42 -188 -37 -186
rect -35 -188 -29 -186
rect -42 -189 -29 -188
rect -65 -205 -63 -203
rect -65 -209 -61 -205
rect -33 -198 -29 -189
rect -65 -211 -64 -209
rect -62 -211 -61 -209
rect -65 -214 -61 -211
rect -164 -221 -163 -219
rect -161 -221 -160 -219
rect -164 -222 -160 -221
rect -50 -216 -44 -209
rect -50 -218 -37 -216
rect -50 -220 -46 -218
rect -44 -220 -37 -218
rect -50 -222 -37 -220
rect -69 -228 -25 -227
rect -69 -230 -62 -228
rect -60 -230 -48 -228
rect -46 -230 -34 -228
rect -32 -230 -25 -228
rect -13 -230 -9 -92
rect 3 -93 10 -92
rect 12 -93 18 -91
rect 20 -93 90 -91
rect 92 -93 98 -91
rect 100 -93 170 -91
rect 172 -93 178 -91
rect 180 -93 250 -91
rect 252 -93 258 -91
rect 260 -93 327 -91
rect 3 -94 327 -93
rect 7 -116 12 -114
rect 7 -118 9 -116
rect 11 -118 12 -116
rect 7 -120 12 -118
rect 7 -131 11 -120
rect 7 -137 19 -131
rect 7 -142 13 -137
rect 7 -144 9 -142
rect 11 -144 13 -142
rect 7 -145 13 -144
rect 63 -117 68 -115
rect 63 -119 65 -117
rect 67 -119 68 -117
rect 63 -121 68 -119
rect 63 -132 67 -121
rect 54 -136 67 -132
rect 71 -127 75 -125
rect 71 -129 72 -127
rect 74 -129 75 -127
rect 71 -140 75 -129
rect 87 -116 92 -114
rect 87 -118 89 -116
rect 91 -118 92 -116
rect 87 -120 92 -118
rect 87 -131 91 -120
rect 87 -137 99 -131
rect 62 -144 75 -140
rect 87 -142 93 -137
rect 87 -144 89 -142
rect 91 -144 93 -142
rect 87 -145 93 -144
rect 143 -117 148 -115
rect 143 -119 145 -117
rect 147 -119 148 -117
rect 143 -121 148 -119
rect 143 -132 147 -121
rect 134 -136 147 -132
rect 151 -127 155 -125
rect 151 -129 152 -127
rect 154 -129 155 -127
rect 151 -140 155 -129
rect 167 -116 172 -114
rect 167 -118 169 -116
rect 171 -118 172 -116
rect 167 -120 172 -118
rect 167 -131 171 -120
rect 167 -137 179 -131
rect 142 -144 155 -140
rect 167 -142 173 -137
rect 167 -144 169 -142
rect 171 -144 173 -142
rect 167 -145 173 -144
rect 223 -117 228 -115
rect 223 -119 225 -117
rect 227 -119 228 -117
rect 223 -121 228 -119
rect 223 -132 227 -121
rect 214 -136 227 -132
rect 231 -127 235 -125
rect 231 -129 232 -127
rect 234 -129 235 -127
rect 231 -140 235 -129
rect 247 -116 252 -114
rect 247 -118 249 -116
rect 251 -118 252 -116
rect 247 -120 252 -118
rect 247 -131 251 -120
rect 247 -137 259 -131
rect 222 -144 235 -140
rect 247 -142 253 -137
rect 247 -144 249 -142
rect 251 -144 253 -142
rect 247 -145 253 -144
rect 303 -117 308 -115
rect 303 -119 305 -117
rect 307 -119 308 -117
rect 303 -121 308 -119
rect 303 -132 307 -121
rect 294 -136 307 -132
rect 311 -127 315 -125
rect 311 -129 312 -127
rect 314 -129 315 -127
rect 311 -140 315 -129
rect 302 -144 315 -140
rect 3 -151 327 -150
rect 341 -151 346 8
rect 3 -153 30 -151
rect 32 -153 70 -151
rect 72 -153 110 -151
rect 112 -153 150 -151
rect 152 -153 190 -151
rect 192 -153 230 -151
rect 232 -153 270 -151
rect 272 -153 310 -151
rect 312 -153 346 -151
rect 3 -155 346 -153
rect 3 -158 327 -155
rect 55 -164 60 -158
rect 3 -165 327 -164
rect 3 -167 4 -165
rect 6 -167 327 -165
rect 3 -169 327 -167
rect 3 -171 30 -169
rect 32 -171 70 -169
rect 72 -171 110 -169
rect 112 -171 150 -169
rect 152 -171 190 -169
rect 192 -171 230 -169
rect 232 -171 270 -169
rect 272 -171 310 -169
rect 312 -171 327 -169
rect 3 -172 327 -171
rect 7 -178 13 -177
rect 7 -180 9 -178
rect 11 -180 13 -178
rect 7 -185 13 -180
rect 7 -191 19 -185
rect 7 -202 11 -191
rect 87 -178 93 -177
rect 62 -182 75 -178
rect 87 -180 89 -178
rect 91 -180 93 -178
rect 54 -190 67 -186
rect 7 -204 12 -202
rect 7 -206 9 -204
rect 11 -206 12 -204
rect 7 -208 12 -206
rect 63 -201 67 -190
rect 71 -193 75 -182
rect 71 -195 72 -193
rect 74 -195 75 -193
rect 71 -197 75 -195
rect 63 -203 68 -201
rect 63 -205 65 -203
rect 67 -205 68 -203
rect 63 -207 68 -205
rect 87 -185 93 -180
rect 87 -191 99 -185
rect 87 -202 91 -191
rect 167 -178 173 -177
rect 142 -182 155 -178
rect 167 -180 169 -178
rect 171 -180 173 -178
rect 134 -190 147 -186
rect 87 -204 92 -202
rect 87 -206 89 -204
rect 91 -206 92 -204
rect 87 -208 92 -206
rect 143 -201 147 -190
rect 151 -193 155 -182
rect 151 -195 152 -193
rect 154 -195 155 -193
rect 151 -197 155 -195
rect 143 -203 148 -201
rect 143 -205 145 -203
rect 147 -205 148 -203
rect 143 -207 148 -205
rect 167 -185 173 -180
rect 167 -191 179 -185
rect 167 -202 171 -191
rect 247 -178 253 -177
rect 222 -182 235 -178
rect 247 -180 249 -178
rect 251 -180 253 -178
rect 214 -190 227 -186
rect 167 -204 172 -202
rect 167 -206 169 -204
rect 171 -206 172 -204
rect 167 -208 172 -206
rect 223 -201 227 -190
rect 231 -193 235 -182
rect 231 -195 232 -193
rect 234 -195 235 -193
rect 231 -197 235 -195
rect 223 -203 228 -201
rect 223 -205 225 -203
rect 227 -205 228 -203
rect 223 -207 228 -205
rect 247 -185 253 -180
rect 247 -191 259 -185
rect 247 -202 251 -191
rect 302 -182 315 -178
rect 294 -190 307 -186
rect 247 -204 252 -202
rect 247 -206 249 -204
rect 251 -206 252 -204
rect 247 -208 252 -206
rect 303 -201 307 -190
rect 311 -193 315 -182
rect 311 -195 312 -193
rect 314 -195 315 -193
rect 311 -197 315 -195
rect 303 -203 308 -201
rect 303 -205 305 -203
rect 307 -205 308 -203
rect 303 -207 308 -205
rect 3 -229 327 -228
rect 3 -230 10 -229
rect -69 -231 10 -230
rect 12 -231 18 -229
rect 20 -231 90 -229
rect 92 -231 98 -229
rect 100 -231 170 -229
rect 172 -231 178 -229
rect 180 -231 250 -229
rect 252 -231 258 -229
rect 260 -231 327 -229
rect -69 -234 327 -231
rect -69 -235 -25 -234
rect 3 -236 327 -234
<< alu2 >>
rect -67 38 -27 39
rect -102 37 -98 38
rect -102 35 -101 37
rect -99 35 -98 37
rect -67 36 -66 38
rect -64 36 321 38
rect -67 35 72 36
rect -102 -94 -98 35
rect -31 34 72 35
rect 74 34 154 36
rect 156 34 235 36
rect 237 34 318 36
rect 320 34 321 36
rect -31 33 321 34
rect -81 30 -35 31
rect -81 29 -39 30
rect -81 27 -80 29
rect -78 28 -39 29
rect -37 28 -35 30
rect -78 27 -35 28
rect -81 26 -35 27
rect -30 10 7 11
rect -92 9 -88 10
rect -92 7 -91 9
rect -89 7 -88 9
rect -30 8 -29 10
rect -27 8 4 10
rect 6 8 7 10
rect -30 7 7 8
rect -92 -2 -88 7
rect -92 -3 -67 -2
rect -92 -5 -70 -3
rect -68 -5 -67 -3
rect -92 -6 -67 -5
rect -93 -18 -89 -17
rect -93 -20 -92 -18
rect -90 -20 -89 -18
rect -93 -55 -89 -20
rect -81 -25 -34 -23
rect -81 -27 -80 -25
rect -78 -27 -38 -25
rect -36 -27 -34 -25
rect -81 -28 -34 -27
rect -66 -33 318 -32
rect -66 -34 72 -33
rect -66 -36 -65 -34
rect -63 -35 72 -34
rect 74 -35 152 -33
rect 154 -35 235 -33
rect 237 -35 315 -33
rect 317 -35 318 -33
rect -63 -36 318 -35
rect -66 -37 318 -36
rect -93 -57 -43 -55
rect -93 -59 -47 -57
rect -45 -59 -43 -57
rect -93 -61 -43 -59
rect -102 -96 -42 -94
rect -102 -98 -46 -96
rect -44 -98 -42 -96
rect -102 -100 -42 -98
rect -65 -119 -13 -118
rect -65 -121 -64 -119
rect -62 -121 -13 -119
rect -65 -122 -13 -121
rect -17 -125 -13 -122
rect -17 -127 315 -125
rect -152 -128 -33 -127
rect -152 -129 -37 -128
rect -152 -131 -151 -129
rect -149 -130 -37 -129
rect -35 -130 -33 -128
rect -149 -131 -33 -130
rect -17 -129 72 -127
rect 74 -129 152 -127
rect 154 -129 232 -127
rect 234 -129 312 -127
rect 314 -129 315 -127
rect -17 -131 315 -129
rect -152 -132 -33 -131
rect -28 -165 7 -164
rect -28 -167 -27 -165
rect -25 -167 4 -165
rect 6 -167 7 -165
rect -28 -168 7 -167
rect -152 -186 -33 -184
rect -152 -188 -151 -186
rect -149 -188 -37 -186
rect -35 -188 -33 -186
rect -152 -189 -33 -188
rect -19 -193 315 -191
rect -19 -195 72 -193
rect 74 -195 152 -193
rect 154 -195 232 -193
rect 234 -195 312 -193
rect 314 -195 315 -193
rect -19 -196 315 -195
rect -20 -197 315 -196
rect -20 -206 -15 -197
rect -65 -209 -15 -206
rect -65 -211 -64 -209
rect -62 -211 -15 -209
rect -65 -212 -15 -211
rect -164 -218 -42 -216
rect -164 -219 -46 -218
rect -164 -221 -163 -219
rect -161 -220 -46 -219
rect -44 -220 -42 -218
rect -161 -221 -42 -220
rect -164 -222 -42 -221
<< ptie >>
rect -128 10 -114 15
rect -128 8 -126 10
rect -124 8 -118 10
rect -116 8 -114 10
rect -66 12 -60 14
rect -66 10 -64 12
rect -62 10 -60 12
rect -66 8 -60 10
rect 28 12 34 14
rect 28 10 30 12
rect 32 10 34 12
rect 28 8 34 10
rect 110 12 116 14
rect 110 10 112 12
rect 114 10 116 12
rect 110 8 116 10
rect 191 12 197 14
rect 191 10 193 12
rect 195 10 197 12
rect 191 8 197 10
rect 274 12 280 14
rect 274 10 276 12
rect 278 10 280 12
rect 274 8 280 10
rect -128 6 -114 8
rect -65 -7 -59 -5
rect -128 -9 -114 -7
rect -128 -11 -126 -9
rect -124 -11 -118 -9
rect -116 -11 -114 -9
rect -65 -9 -63 -7
rect -61 -9 -59 -7
rect -65 -11 -59 -9
rect 28 -9 34 -7
rect -128 -16 -114 -11
rect 28 -11 30 -9
rect 32 -11 34 -9
rect 28 -13 34 -11
rect 108 -9 114 -7
rect 108 -11 110 -9
rect 112 -11 114 -9
rect 108 -13 114 -11
rect 191 -9 197 -7
rect 191 -11 193 -9
rect 195 -11 197 -9
rect 191 -13 197 -11
rect 271 -9 277 -7
rect 271 -11 273 -9
rect 275 -11 277 -9
rect 271 -13 277 -11
rect -64 -146 -58 -144
rect -64 -148 -62 -146
rect -60 -148 -58 -146
rect -64 -150 -58 -148
rect 28 -151 34 -149
rect 28 -153 30 -151
rect 32 -153 34 -151
rect 28 -155 34 -153
rect 108 -151 114 -149
rect 108 -153 110 -151
rect 112 -153 114 -151
rect 108 -155 114 -153
rect 188 -151 194 -149
rect 188 -153 190 -151
rect 192 -153 194 -151
rect 188 -155 194 -153
rect 268 -151 274 -149
rect 268 -153 270 -151
rect 272 -153 274 -151
rect 268 -155 274 -153
rect -64 -168 -58 -166
rect -64 -170 -62 -168
rect -60 -170 -58 -168
rect -64 -172 -58 -170
rect 28 -169 34 -167
rect 28 -171 30 -169
rect 32 -171 34 -169
rect 28 -173 34 -171
rect 108 -169 114 -167
rect 108 -171 110 -169
rect 112 -171 114 -169
rect 108 -173 114 -171
rect 188 -169 194 -167
rect 188 -171 190 -169
rect 192 -171 194 -169
rect 188 -173 194 -171
rect 268 -169 274 -167
rect 268 -171 270 -169
rect 272 -171 274 -169
rect 268 -173 274 -171
<< ntie >>
rect -66 72 -32 74
rect -119 70 -113 72
rect -119 68 -117 70
rect -115 68 -113 70
rect -66 70 -64 72
rect -62 70 -50 72
rect -48 70 -36 72
rect -34 70 -32 72
rect -66 68 -32 70
rect 8 72 22 74
rect 8 70 10 72
rect 12 70 18 72
rect 20 70 22 72
rect 8 68 22 70
rect -119 65 -113 68
rect 90 72 104 74
rect 90 70 92 72
rect 94 70 100 72
rect 102 70 104 72
rect 90 68 104 70
rect 171 72 185 74
rect 171 70 173 72
rect 175 70 181 72
rect 183 70 185 72
rect 171 68 185 70
rect 254 72 268 74
rect 254 70 256 72
rect 258 70 264 72
rect 266 70 268 72
rect 254 68 268 70
rect -119 -69 -113 -66
rect -119 -71 -117 -69
rect -115 -71 -113 -69
rect -65 -67 -31 -65
rect -65 -69 -63 -67
rect -61 -69 -49 -67
rect -47 -69 -35 -67
rect -33 -69 -31 -67
rect -65 -71 -31 -69
rect 8 -69 22 -67
rect 8 -71 10 -69
rect 12 -71 18 -69
rect 20 -71 22 -69
rect -119 -73 -113 -71
rect 8 -73 22 -71
rect 88 -69 102 -67
rect 88 -71 90 -69
rect 92 -71 98 -69
rect 100 -71 102 -69
rect 88 -73 102 -71
rect 171 -69 185 -67
rect 171 -71 173 -69
rect 175 -71 181 -69
rect 183 -71 185 -69
rect 171 -73 185 -71
rect 251 -69 265 -67
rect 251 -71 253 -69
rect 255 -71 261 -69
rect 263 -71 265 -69
rect 251 -73 265 -71
rect -64 -86 -30 -84
rect -64 -88 -62 -86
rect -60 -88 -48 -86
rect -46 -88 -34 -86
rect -32 -88 -30 -86
rect -64 -90 -30 -88
rect 8 -91 22 -89
rect 8 -93 10 -91
rect 12 -93 18 -91
rect 20 -93 22 -91
rect 8 -95 22 -93
rect 88 -91 102 -89
rect 88 -93 90 -91
rect 92 -93 98 -91
rect 100 -93 102 -91
rect 88 -95 102 -93
rect 168 -91 182 -89
rect 168 -93 170 -91
rect 172 -93 178 -91
rect 180 -93 182 -91
rect 168 -95 182 -93
rect 248 -91 262 -89
rect 248 -93 250 -91
rect 252 -93 258 -91
rect 260 -93 262 -91
rect 248 -95 262 -93
rect -64 -228 -30 -226
rect -64 -230 -62 -228
rect -60 -230 -48 -228
rect -46 -230 -34 -228
rect -32 -230 -30 -228
rect -64 -232 -30 -230
rect 8 -229 22 -227
rect 8 -231 10 -229
rect 12 -231 18 -229
rect 20 -231 22 -229
rect 8 -233 22 -231
rect 88 -229 102 -227
rect 88 -231 90 -229
rect 92 -231 98 -229
rect 100 -231 102 -229
rect 88 -233 102 -231
rect 168 -229 182 -227
rect 168 -231 170 -229
rect 172 -231 178 -229
rect 180 -231 182 -229
rect 168 -233 182 -231
rect 248 -229 262 -227
rect 248 -231 250 -229
rect 252 -231 258 -229
rect 260 -231 262 -229
rect 248 -233 262 -231
<< nmos >>
rect -122 23 -120 29
rect -60 20 -58 26
rect -48 14 -46 23
rect -41 14 -39 23
rect 29 25 31 31
rect 15 15 17 21
rect 40 19 42 25
rect 47 19 49 25
rect 57 19 59 25
rect 64 19 66 25
rect 74 23 76 29
rect 111 25 113 31
rect 97 15 99 21
rect 122 19 124 25
rect 129 19 131 25
rect 139 19 141 25
rect 146 19 148 25
rect 156 23 158 29
rect 192 25 194 31
rect 178 15 180 21
rect 203 19 205 25
rect 210 19 212 25
rect 220 19 222 25
rect 227 19 229 25
rect 237 23 239 29
rect 275 25 277 31
rect 261 15 263 21
rect 286 19 288 25
rect 293 19 295 25
rect 303 19 305 25
rect 310 19 312 25
rect 320 23 322 29
rect -59 -23 -57 -17
rect -47 -20 -45 -11
rect -40 -20 -38 -11
rect 15 -20 17 -14
rect -122 -30 -120 -24
rect 40 -24 42 -18
rect 47 -24 49 -18
rect 57 -24 59 -18
rect 64 -24 66 -18
rect 95 -20 97 -14
rect 29 -30 31 -24
rect 74 -28 76 -22
rect 120 -24 122 -18
rect 127 -24 129 -18
rect 137 -24 139 -18
rect 144 -24 146 -18
rect 178 -20 180 -14
rect 109 -30 111 -24
rect 154 -28 156 -22
rect 203 -24 205 -18
rect 210 -24 212 -18
rect 220 -24 222 -18
rect 227 -24 229 -18
rect 258 -20 260 -14
rect 192 -30 194 -24
rect 237 -28 239 -22
rect 283 -24 285 -18
rect 290 -24 292 -18
rect 300 -24 302 -18
rect 307 -24 309 -18
rect 272 -30 274 -24
rect 317 -28 319 -22
rect -58 -138 -56 -132
rect -46 -144 -44 -135
rect -39 -144 -37 -135
rect 29 -138 31 -132
rect 15 -148 17 -142
rect 40 -144 42 -138
rect 47 -144 49 -138
rect 57 -144 59 -138
rect 64 -144 66 -138
rect 74 -140 76 -134
rect 109 -138 111 -132
rect 95 -148 97 -142
rect 120 -144 122 -138
rect 127 -144 129 -138
rect 137 -144 139 -138
rect 144 -144 146 -138
rect 154 -140 156 -134
rect 189 -138 191 -132
rect 175 -148 177 -142
rect 200 -144 202 -138
rect 207 -144 209 -138
rect 217 -144 219 -138
rect 224 -144 226 -138
rect 234 -140 236 -134
rect 269 -138 271 -132
rect 255 -148 257 -142
rect 280 -144 282 -138
rect 287 -144 289 -138
rect 297 -144 299 -138
rect 304 -144 306 -138
rect 314 -140 316 -134
rect -58 -184 -56 -178
rect -46 -181 -44 -172
rect -39 -181 -37 -172
rect 15 -180 17 -174
rect 40 -184 42 -178
rect 47 -184 49 -178
rect 57 -184 59 -178
rect 64 -184 66 -178
rect 95 -180 97 -174
rect 29 -190 31 -184
rect 74 -188 76 -182
rect 120 -184 122 -178
rect 127 -184 129 -178
rect 137 -184 139 -178
rect 144 -184 146 -178
rect 175 -180 177 -174
rect 109 -190 111 -184
rect 154 -188 156 -182
rect 200 -184 202 -178
rect 207 -184 209 -178
rect 217 -184 219 -178
rect 224 -184 226 -178
rect 255 -180 257 -174
rect 189 -190 191 -184
rect 234 -188 236 -182
rect 280 -184 282 -178
rect 287 -184 289 -178
rect 297 -184 299 -178
rect 304 -184 306 -178
rect 269 -190 271 -184
rect 314 -188 316 -182
<< pmos >>
rect -122 41 -120 53
rect -60 43 -58 55
rect 40 59 42 65
rect 47 59 49 65
rect -50 43 -48 53
rect -40 43 -38 53
rect 14 43 16 55
rect 24 43 26 55
rect 57 53 59 65
rect 64 53 66 65
rect 74 53 76 65
rect 122 59 124 65
rect 129 59 131 65
rect 96 43 98 55
rect 106 43 108 55
rect 139 53 141 65
rect 146 53 148 65
rect 156 53 158 65
rect 203 59 205 65
rect 210 59 212 65
rect 177 43 179 55
rect 187 43 189 55
rect 220 53 222 65
rect 227 53 229 65
rect 237 53 239 65
rect 286 59 288 65
rect 293 59 295 65
rect 260 43 262 55
rect 270 43 272 55
rect 303 53 305 65
rect 310 53 312 65
rect 320 53 322 65
rect -122 -54 -120 -42
rect -59 -52 -57 -40
rect -49 -50 -47 -40
rect -39 -50 -37 -40
rect 14 -54 16 -42
rect 24 -54 26 -42
rect 40 -64 42 -58
rect 47 -64 49 -58
rect 57 -64 59 -52
rect 64 -64 66 -52
rect 74 -64 76 -52
rect 94 -54 96 -42
rect 104 -54 106 -42
rect 120 -64 122 -58
rect 127 -64 129 -58
rect 137 -64 139 -52
rect 144 -64 146 -52
rect 154 -64 156 -52
rect 177 -54 179 -42
rect 187 -54 189 -42
rect 203 -64 205 -58
rect 210 -64 212 -58
rect 220 -64 222 -52
rect 227 -64 229 -52
rect 237 -64 239 -52
rect 257 -54 259 -42
rect 267 -54 269 -42
rect 283 -64 285 -58
rect 290 -64 292 -58
rect 300 -64 302 -52
rect 307 -64 309 -52
rect 317 -64 319 -52
rect -58 -115 -56 -103
rect -48 -115 -46 -105
rect -38 -115 -36 -105
rect 40 -104 42 -98
rect 47 -104 49 -98
rect 14 -120 16 -108
rect 24 -120 26 -108
rect 57 -110 59 -98
rect 64 -110 66 -98
rect 74 -110 76 -98
rect 120 -104 122 -98
rect 127 -104 129 -98
rect 94 -120 96 -108
rect 104 -120 106 -108
rect 137 -110 139 -98
rect 144 -110 146 -98
rect 154 -110 156 -98
rect 200 -104 202 -98
rect 207 -104 209 -98
rect 174 -120 176 -108
rect 184 -120 186 -108
rect 217 -110 219 -98
rect 224 -110 226 -98
rect 234 -110 236 -98
rect 280 -104 282 -98
rect 287 -104 289 -98
rect 254 -120 256 -108
rect 264 -120 266 -108
rect 297 -110 299 -98
rect 304 -110 306 -98
rect 314 -110 316 -98
rect -58 -213 -56 -201
rect -48 -211 -46 -201
rect -38 -211 -36 -201
rect 14 -214 16 -202
rect 24 -214 26 -202
rect 40 -224 42 -218
rect 47 -224 49 -218
rect 57 -224 59 -212
rect 64 -224 66 -212
rect 74 -224 76 -212
rect 94 -214 96 -202
rect 104 -214 106 -202
rect 120 -224 122 -218
rect 127 -224 129 -218
rect 137 -224 139 -212
rect 144 -224 146 -212
rect 154 -224 156 -212
rect 174 -214 176 -202
rect 184 -214 186 -202
rect 200 -224 202 -218
rect 207 -224 209 -218
rect 217 -224 219 -212
rect 224 -224 226 -212
rect 234 -224 236 -212
rect 254 -214 256 -202
rect 264 -214 266 -202
rect 280 -224 282 -218
rect 287 -224 289 -218
rect 297 -224 299 -212
rect 304 -224 306 -212
rect 314 -224 316 -212
<< polyct0 >>
rect 38 52 40 54
rect -58 36 -56 38
rect 32 36 34 38
rect 55 46 57 48
rect 48 30 50 32
rect 120 52 122 54
rect 114 36 116 38
rect 137 46 139 48
rect 130 30 132 32
rect 201 52 203 54
rect 195 36 197 38
rect 218 46 220 48
rect 211 30 213 32
rect 284 52 286 54
rect 278 36 280 38
rect 301 46 303 48
rect 294 30 296 32
rect -57 -35 -55 -33
rect 32 -37 34 -35
rect 48 -31 50 -29
rect 38 -53 40 -51
rect 112 -37 114 -35
rect 55 -47 57 -45
rect 128 -31 130 -29
rect 118 -53 120 -51
rect 195 -37 197 -35
rect 135 -47 137 -45
rect 211 -31 213 -29
rect 201 -53 203 -51
rect 275 -37 277 -35
rect 218 -47 220 -45
rect 291 -31 293 -29
rect 281 -53 283 -51
rect 298 -47 300 -45
rect -56 -122 -54 -120
rect 38 -111 40 -109
rect 32 -127 34 -125
rect 55 -117 57 -115
rect 48 -133 50 -131
rect 118 -111 120 -109
rect 112 -127 114 -125
rect 135 -117 137 -115
rect 128 -133 130 -131
rect 198 -111 200 -109
rect 192 -127 194 -125
rect 215 -117 217 -115
rect 208 -133 210 -131
rect 278 -111 280 -109
rect 272 -127 274 -125
rect 295 -117 297 -115
rect 288 -133 290 -131
rect -56 -196 -54 -194
rect 32 -197 34 -195
rect 48 -191 50 -189
rect 38 -213 40 -211
rect 112 -197 114 -195
rect 55 -207 57 -205
rect 128 -191 130 -189
rect 118 -213 120 -211
rect 192 -197 194 -195
rect 135 -207 137 -205
rect 208 -191 210 -189
rect 198 -213 200 -211
rect 272 -197 274 -195
rect 215 -207 217 -205
rect 288 -191 290 -189
rect 278 -213 280 -211
rect 295 -207 297 -205
<< polyct1 >>
rect -48 60 -46 62
rect -120 58 -118 60
rect -39 28 -37 30
rect 65 44 67 46
rect 72 34 74 36
rect 147 44 149 46
rect 154 34 156 36
rect 228 44 230 46
rect 235 34 237 36
rect 311 44 313 46
rect 318 34 320 36
rect -38 -27 -36 -25
rect -120 -61 -118 -59
rect -47 -59 -45 -57
rect 72 -35 74 -33
rect 65 -45 67 -43
rect 152 -35 154 -33
rect 145 -45 147 -43
rect 235 -35 237 -33
rect 228 -45 230 -43
rect 315 -35 317 -33
rect 308 -45 310 -43
rect -46 -98 -44 -96
rect -37 -130 -35 -128
rect 65 -119 67 -117
rect 72 -129 74 -127
rect 145 -119 147 -117
rect 152 -129 154 -127
rect 225 -119 227 -117
rect 232 -129 234 -127
rect 305 -119 307 -117
rect 312 -129 314 -127
rect -37 -188 -35 -186
rect -46 -220 -44 -218
rect 72 -195 74 -193
rect 65 -205 67 -203
rect 152 -195 154 -193
rect 145 -205 147 -203
rect 232 -195 234 -193
rect 225 -205 227 -203
rect 312 -195 314 -193
rect 305 -205 307 -203
<< ndifct0 >>
rect -117 25 -115 27
rect -36 19 -34 21
rect 24 27 26 29
rect 34 27 36 29
rect 52 21 54 23
rect 79 25 81 27
rect 20 17 22 19
rect 106 27 108 29
rect 116 27 118 29
rect 134 21 136 23
rect 161 25 163 27
rect 102 17 104 19
rect 187 27 189 29
rect 197 27 199 29
rect 215 21 217 23
rect 242 25 244 27
rect 183 17 185 19
rect 270 27 272 29
rect 280 27 282 29
rect 298 21 300 23
rect 325 25 327 27
rect 266 17 268 19
rect -35 -18 -33 -16
rect 20 -18 22 -16
rect -117 -28 -115 -26
rect 52 -22 54 -20
rect 100 -18 102 -16
rect 24 -28 26 -26
rect 34 -28 36 -26
rect 79 -26 81 -24
rect 132 -22 134 -20
rect 183 -18 185 -16
rect 104 -28 106 -26
rect 114 -28 116 -26
rect 159 -26 161 -24
rect 215 -22 217 -20
rect 263 -18 265 -16
rect 187 -28 189 -26
rect 197 -28 199 -26
rect 242 -26 244 -24
rect 295 -22 297 -20
rect 267 -28 269 -26
rect 277 -28 279 -26
rect 322 -26 324 -24
rect -34 -139 -32 -137
rect 24 -136 26 -134
rect 34 -136 36 -134
rect 52 -142 54 -140
rect 79 -138 81 -136
rect 20 -146 22 -144
rect 104 -136 106 -134
rect 114 -136 116 -134
rect 132 -142 134 -140
rect 159 -138 161 -136
rect 100 -146 102 -144
rect 184 -136 186 -134
rect 194 -136 196 -134
rect 212 -142 214 -140
rect 239 -138 241 -136
rect 180 -146 182 -144
rect 264 -136 266 -134
rect 274 -136 276 -134
rect 292 -142 294 -140
rect 319 -138 321 -136
rect 260 -146 262 -144
rect -34 -179 -32 -177
rect 20 -178 22 -176
rect 52 -182 54 -180
rect 100 -178 102 -176
rect 24 -188 26 -186
rect 34 -188 36 -186
rect 79 -186 81 -184
rect 132 -182 134 -180
rect 180 -178 182 -176
rect 104 -188 106 -186
rect 114 -188 116 -186
rect 159 -186 161 -184
rect 212 -182 214 -180
rect 260 -178 262 -176
rect 184 -188 186 -186
rect 194 -188 196 -186
rect 239 -186 241 -184
rect 292 -182 294 -180
rect 264 -188 266 -186
rect 274 -188 276 -186
rect 319 -186 321 -184
<< ndifct1 >>
rect -127 25 -125 27
rect -65 22 -63 24
rect 9 19 11 21
rect -54 10 -52 12
rect 91 19 93 21
rect 70 10 72 12
rect 172 19 174 21
rect 152 10 154 12
rect 255 19 257 21
rect 233 10 235 12
rect 316 10 318 12
rect -53 -9 -51 -7
rect -64 -21 -62 -19
rect 70 -11 72 -9
rect 9 -20 11 -18
rect 150 -11 152 -9
rect -127 -28 -125 -26
rect 89 -20 91 -18
rect 233 -11 235 -9
rect 172 -20 174 -18
rect 313 -11 315 -9
rect 252 -20 254 -18
rect -63 -136 -61 -134
rect 9 -144 11 -142
rect -52 -148 -50 -146
rect 89 -144 91 -142
rect 70 -153 72 -151
rect 169 -144 171 -142
rect 150 -153 152 -151
rect 249 -144 251 -142
rect 230 -153 232 -151
rect 310 -153 312 -151
rect -52 -170 -50 -168
rect -63 -182 -61 -180
rect 70 -171 72 -169
rect 9 -180 11 -178
rect 150 -171 152 -169
rect 89 -180 91 -178
rect 230 -171 232 -169
rect 169 -180 171 -178
rect 310 -171 312 -169
rect 249 -180 251 -178
<< ntiect1 >>
rect -117 68 -115 70
rect -64 70 -62 72
rect -50 70 -48 72
rect -36 70 -34 72
rect 10 70 12 72
rect 18 70 20 72
rect 92 70 94 72
rect 100 70 102 72
rect 173 70 175 72
rect 181 70 183 72
rect 256 70 258 72
rect 264 70 266 72
rect -117 -71 -115 -69
rect -63 -69 -61 -67
rect -49 -69 -47 -67
rect -35 -69 -33 -67
rect 10 -71 12 -69
rect 18 -71 20 -69
rect 90 -71 92 -69
rect 98 -71 100 -69
rect 173 -71 175 -69
rect 181 -71 183 -69
rect 253 -71 255 -69
rect 261 -71 263 -69
rect -62 -88 -60 -86
rect -48 -88 -46 -86
rect -34 -88 -32 -86
rect 10 -93 12 -91
rect 18 -93 20 -91
rect 90 -93 92 -91
rect 98 -93 100 -91
rect 170 -93 172 -91
rect 178 -93 180 -91
rect 250 -93 252 -91
rect 258 -93 260 -91
rect -62 -230 -60 -228
rect -48 -230 -46 -228
rect -34 -230 -32 -228
rect 10 -231 12 -229
rect 18 -231 20 -229
rect 90 -231 92 -229
rect 98 -231 100 -229
rect 170 -231 172 -229
rect 178 -231 180 -229
rect 250 -231 252 -229
rect 258 -231 260 -229
<< ptiect1 >>
rect -126 8 -124 10
rect -118 8 -116 10
rect -64 10 -62 12
rect 30 10 32 12
rect 112 10 114 12
rect 193 10 195 12
rect 276 10 278 12
rect -126 -11 -124 -9
rect -118 -11 -116 -9
rect -63 -9 -61 -7
rect 30 -11 32 -9
rect 110 -11 112 -9
rect 193 -11 195 -9
rect 273 -11 275 -9
rect -62 -148 -60 -146
rect 30 -153 32 -151
rect 110 -153 112 -151
rect 190 -153 192 -151
rect 270 -153 272 -151
rect -62 -170 -60 -168
rect 30 -171 32 -169
rect 110 -171 112 -169
rect 190 -171 192 -169
rect 270 -171 272 -169
<< pdifct0 >>
rect 35 61 37 63
rect 52 61 54 63
rect -55 45 -53 47
rect -45 45 -43 47
rect -35 49 -33 51
rect 19 51 21 53
rect 29 51 31 53
rect 69 61 71 63
rect 117 61 119 63
rect 79 55 81 57
rect 134 61 136 63
rect 101 51 103 53
rect 111 51 113 53
rect 151 61 153 63
rect 198 61 200 63
rect 161 55 163 57
rect 215 61 217 63
rect 182 51 184 53
rect 192 51 194 53
rect 232 61 234 63
rect 281 61 283 63
rect 242 55 244 57
rect 298 61 300 63
rect 265 51 267 53
rect 275 51 277 53
rect 315 61 317 63
rect 325 55 327 57
rect -54 -44 -52 -42
rect -44 -44 -42 -42
rect -34 -48 -32 -46
rect 19 -52 21 -50
rect 29 -52 31 -50
rect 35 -62 37 -60
rect 52 -62 54 -60
rect 69 -62 71 -60
rect 99 -52 101 -50
rect 109 -52 111 -50
rect 79 -56 81 -54
rect 115 -62 117 -60
rect 132 -62 134 -60
rect 149 -62 151 -60
rect 182 -52 184 -50
rect 192 -52 194 -50
rect 159 -56 161 -54
rect 198 -62 200 -60
rect 215 -62 217 -60
rect 232 -62 234 -60
rect 262 -52 264 -50
rect 272 -52 274 -50
rect 242 -56 244 -54
rect 278 -62 280 -60
rect 295 -62 297 -60
rect 312 -62 314 -60
rect 322 -56 324 -54
rect 35 -102 37 -100
rect -53 -113 -51 -111
rect -43 -113 -41 -111
rect -33 -109 -31 -107
rect 52 -102 54 -100
rect 19 -112 21 -110
rect 29 -112 31 -110
rect 69 -102 71 -100
rect 115 -102 117 -100
rect 79 -108 81 -106
rect 132 -102 134 -100
rect 99 -112 101 -110
rect 109 -112 111 -110
rect 149 -102 151 -100
rect 195 -102 197 -100
rect 159 -108 161 -106
rect 212 -102 214 -100
rect 179 -112 181 -110
rect 189 -112 191 -110
rect 229 -102 231 -100
rect 275 -102 277 -100
rect 239 -108 241 -106
rect 292 -102 294 -100
rect 259 -112 261 -110
rect 269 -112 271 -110
rect 309 -102 311 -100
rect 319 -108 321 -106
rect -53 -205 -51 -203
rect -43 -205 -41 -203
rect -33 -209 -31 -207
rect 19 -212 21 -210
rect 29 -212 31 -210
rect 35 -222 37 -220
rect 52 -222 54 -220
rect 69 -222 71 -220
rect 99 -212 101 -210
rect 109 -212 111 -210
rect 79 -216 81 -214
rect 115 -222 117 -220
rect 132 -222 134 -220
rect 149 -222 151 -220
rect 179 -212 181 -210
rect 189 -212 191 -210
rect 159 -216 161 -214
rect 195 -222 197 -220
rect 212 -222 214 -220
rect 229 -222 231 -220
rect 259 -212 261 -210
rect 269 -212 271 -210
rect 239 -216 241 -214
rect 275 -222 277 -220
rect 292 -222 294 -220
rect 309 -222 311 -220
rect 319 -216 321 -214
<< pdifct1 >>
rect -127 68 -125 70
rect -117 43 -115 45
rect -65 45 -63 47
rect 9 45 11 47
rect 91 45 93 47
rect 172 45 174 47
rect 255 45 257 47
rect -117 -46 -115 -44
rect -64 -44 -62 -42
rect 9 -46 11 -44
rect 89 -46 91 -44
rect 172 -46 174 -44
rect 252 -46 254 -44
rect -127 -71 -125 -69
rect -63 -113 -61 -111
rect 9 -118 11 -116
rect 89 -118 91 -116
rect 169 -118 171 -116
rect 249 -118 251 -116
rect -63 -205 -61 -203
rect 9 -206 11 -204
rect 89 -206 91 -204
rect 169 -206 171 -204
rect 249 -206 251 -204
<< alu0 >>
rect -59 62 -55 69
rect -63 43 -62 49
rect -59 48 -55 60
rect -36 51 -32 69
rect -36 49 -35 51
rect -33 49 -32 51
rect -59 47 -51 48
rect -59 45 -55 47
rect -53 45 -51 47
rect -59 44 -51 45
rect -47 47 -41 48
rect -36 47 -32 49
rect -47 45 -45 47
rect -43 45 -41 47
rect -47 39 -41 45
rect -119 27 -113 28
rect -119 25 -117 27
rect -115 25 -113 27
rect -119 11 -113 25
rect -119 -17 -113 -12
rect -119 -26 -113 -21
rect -119 -28 -117 -26
rect -115 -28 -113 -26
rect -119 -29 -113 -28
rect -60 38 -41 39
rect -60 36 -58 38
rect -56 36 -41 38
rect -60 35 -41 36
rect -63 24 -62 26
rect -51 22 -47 35
rect -51 21 -32 22
rect -51 19 -36 21
rect -34 19 -32 21
rect -51 18 -32 19
rect -50 -16 -31 -15
rect -50 -18 -35 -16
rect -33 -18 -31 -16
rect -50 -19 -31 -18
rect -62 -23 -61 -21
rect -50 -32 -46 -19
rect -59 -33 -40 -32
rect -59 -35 -57 -33
rect -55 -35 -40 -33
rect -59 -36 -40 -35
rect -62 -46 -61 -40
rect -58 -42 -50 -41
rect -58 -44 -54 -42
rect -52 -44 -50 -42
rect -58 -45 -50 -44
rect -46 -42 -40 -36
rect -46 -44 -44 -42
rect -42 -44 -40 -42
rect -46 -45 -40 -44
rect -58 -66 -54 -45
rect -35 -46 -31 -44
rect -35 -48 -34 -46
rect -32 -48 -31 -46
rect -35 -66 -31 -48
rect 17 53 23 69
rect 34 63 38 69
rect 34 61 35 63
rect 37 61 38 63
rect 34 59 38 61
rect 46 63 56 64
rect 46 61 52 63
rect 54 61 56 63
rect 46 60 56 61
rect 68 63 72 69
rect 68 61 69 63
rect 71 61 72 63
rect 17 51 19 53
rect 21 51 23 53
rect 17 50 23 51
rect 28 54 42 55
rect 28 53 38 54
rect 28 51 29 53
rect 31 52 38 53
rect 40 52 42 54
rect 31 51 42 52
rect 28 47 32 51
rect 46 47 50 60
rect 68 59 72 61
rect 78 57 82 59
rect 78 55 79 57
rect 81 55 82 57
rect 23 43 32 47
rect 40 43 50 47
rect 54 51 83 55
rect 54 48 58 51
rect 54 46 55 48
rect 57 46 58 48
rect 23 29 27 43
rect 40 39 44 43
rect 54 39 58 46
rect 30 38 44 39
rect 30 36 32 38
rect 34 36 44 38
rect 30 35 44 36
rect 23 27 24 29
rect 26 27 27 29
rect 23 25 27 27
rect 33 29 37 31
rect 33 27 34 29
rect 36 27 37 29
rect 19 19 23 21
rect 19 17 20 19
rect 22 17 23 19
rect 19 13 23 17
rect 33 13 37 27
rect 40 24 44 35
rect 47 35 58 39
rect 47 32 51 35
rect 47 30 48 32
rect 50 30 51 32
rect 47 28 51 30
rect 40 23 56 24
rect 79 29 83 51
rect 99 53 105 69
rect 116 63 120 69
rect 116 61 117 63
rect 119 61 120 63
rect 116 59 120 61
rect 128 63 138 64
rect 128 61 134 63
rect 136 61 138 63
rect 128 60 138 61
rect 150 63 154 69
rect 150 61 151 63
rect 153 61 154 63
rect 99 51 101 53
rect 103 51 105 53
rect 99 50 105 51
rect 110 54 124 55
rect 110 53 120 54
rect 110 51 111 53
rect 113 52 120 53
rect 122 52 124 54
rect 113 51 124 52
rect 78 27 83 29
rect 78 25 79 27
rect 81 25 83 27
rect 78 23 83 25
rect 110 47 114 51
rect 128 47 132 60
rect 150 59 154 61
rect 160 57 164 59
rect 160 55 161 57
rect 163 55 164 57
rect 105 43 114 47
rect 122 43 132 47
rect 136 51 165 55
rect 136 48 140 51
rect 136 46 137 48
rect 139 46 140 48
rect 105 29 109 43
rect 122 39 126 43
rect 136 39 140 46
rect 112 38 126 39
rect 112 36 114 38
rect 116 36 126 38
rect 112 35 126 36
rect 105 27 106 29
rect 108 27 109 29
rect 40 21 52 23
rect 54 21 56 23
rect 40 20 56 21
rect 105 25 109 27
rect 115 29 119 31
rect 115 27 116 29
rect 118 27 119 29
rect 101 19 105 21
rect 101 17 102 19
rect 104 17 105 19
rect 101 13 105 17
rect 115 13 119 27
rect 122 24 126 35
rect 129 35 140 39
rect 129 32 133 35
rect 129 30 130 32
rect 132 30 133 32
rect 129 28 133 30
rect 122 23 138 24
rect 161 29 165 51
rect 180 53 186 69
rect 197 63 201 69
rect 197 61 198 63
rect 200 61 201 63
rect 197 59 201 61
rect 209 63 219 64
rect 209 61 215 63
rect 217 61 219 63
rect 209 60 219 61
rect 231 63 235 69
rect 231 61 232 63
rect 234 61 235 63
rect 180 51 182 53
rect 184 51 186 53
rect 180 50 186 51
rect 191 54 205 55
rect 191 53 201 54
rect 191 51 192 53
rect 194 52 201 53
rect 203 52 205 54
rect 194 51 205 52
rect 160 27 165 29
rect 160 25 161 27
rect 163 25 165 27
rect 160 23 165 25
rect 191 47 195 51
rect 209 47 213 60
rect 231 59 235 61
rect 241 57 245 59
rect 241 55 242 57
rect 244 55 245 57
rect 186 43 195 47
rect 203 43 213 47
rect 217 51 246 55
rect 217 48 221 51
rect 217 46 218 48
rect 220 46 221 48
rect 186 29 190 43
rect 203 39 207 43
rect 217 39 221 46
rect 193 38 207 39
rect 193 36 195 38
rect 197 36 207 38
rect 193 35 207 36
rect 186 27 187 29
rect 189 27 190 29
rect 122 21 134 23
rect 136 21 138 23
rect 122 20 138 21
rect 186 25 190 27
rect 196 29 200 31
rect 196 27 197 29
rect 199 27 200 29
rect 182 19 186 21
rect 182 17 183 19
rect 185 17 186 19
rect 182 13 186 17
rect 196 13 200 27
rect 203 24 207 35
rect 210 35 221 39
rect 210 32 214 35
rect 210 30 211 32
rect 213 30 214 32
rect 210 28 214 30
rect 203 23 219 24
rect 242 29 246 51
rect 263 53 269 69
rect 280 63 284 69
rect 280 61 281 63
rect 283 61 284 63
rect 280 59 284 61
rect 292 63 302 64
rect 292 61 298 63
rect 300 61 302 63
rect 292 60 302 61
rect 314 63 318 69
rect 314 61 315 63
rect 317 61 318 63
rect 263 51 265 53
rect 267 51 269 53
rect 263 50 269 51
rect 274 54 288 55
rect 274 53 284 54
rect 274 51 275 53
rect 277 52 284 53
rect 286 52 288 54
rect 277 51 288 52
rect 241 27 246 29
rect 241 25 242 27
rect 244 25 246 27
rect 241 23 246 25
rect 274 47 278 51
rect 292 47 296 60
rect 314 59 318 61
rect 324 57 328 59
rect 324 55 325 57
rect 327 55 328 57
rect 269 43 278 47
rect 286 43 296 47
rect 300 51 329 55
rect 300 48 304 51
rect 300 46 301 48
rect 303 46 304 48
rect 269 29 273 43
rect 286 39 290 43
rect 300 39 304 46
rect 276 38 290 39
rect 276 36 278 38
rect 280 36 290 38
rect 276 35 290 36
rect 269 27 270 29
rect 272 27 273 29
rect 203 21 215 23
rect 217 21 219 23
rect 203 20 219 21
rect 269 25 273 27
rect 279 29 283 31
rect 279 27 280 29
rect 282 27 283 29
rect 265 19 269 21
rect 265 17 266 19
rect 268 17 269 19
rect 265 13 269 17
rect 279 13 283 27
rect 286 24 290 35
rect 293 35 304 39
rect 293 32 297 35
rect 293 30 294 32
rect 296 30 297 32
rect 293 28 297 30
rect 286 23 302 24
rect 325 29 329 51
rect 324 27 329 29
rect 324 25 325 27
rect 327 25 329 27
rect 324 23 329 25
rect 286 21 298 23
rect 300 21 302 23
rect 286 20 302 21
rect 19 -16 23 -12
rect 19 -18 20 -16
rect 22 -18 23 -16
rect 19 -20 23 -18
rect 23 -26 27 -24
rect 23 -28 24 -26
rect 26 -28 27 -26
rect 23 -42 27 -28
rect 33 -26 37 -12
rect 99 -16 103 -12
rect 33 -28 34 -26
rect 36 -28 37 -26
rect 33 -30 37 -28
rect 40 -20 56 -19
rect 40 -22 52 -20
rect 54 -22 56 -20
rect 99 -18 100 -16
rect 102 -18 103 -16
rect 99 -20 103 -18
rect 40 -23 56 -22
rect 40 -34 44 -23
rect 30 -35 44 -34
rect 30 -37 32 -35
rect 34 -37 44 -35
rect 30 -38 44 -37
rect 47 -29 51 -27
rect 47 -31 48 -29
rect 50 -31 51 -29
rect 47 -34 51 -31
rect 47 -38 58 -34
rect 40 -42 44 -38
rect 23 -46 32 -42
rect 40 -46 50 -42
rect 17 -50 23 -49
rect 17 -52 19 -50
rect 21 -52 23 -50
rect 17 -68 23 -52
rect 28 -50 32 -46
rect 28 -52 29 -50
rect 31 -51 42 -50
rect 31 -52 38 -51
rect 28 -53 38 -52
rect 40 -53 42 -51
rect 28 -54 42 -53
rect 34 -60 38 -58
rect 34 -62 35 -60
rect 37 -62 38 -60
rect 34 -68 38 -62
rect 46 -59 50 -46
rect 54 -45 58 -38
rect 54 -47 55 -45
rect 57 -47 58 -45
rect 78 -24 83 -22
rect 78 -26 79 -24
rect 81 -26 83 -24
rect 78 -28 83 -26
rect 54 -50 58 -47
rect 79 -50 83 -28
rect 103 -26 107 -24
rect 103 -28 104 -26
rect 106 -28 107 -26
rect 103 -42 107 -28
rect 113 -26 117 -12
rect 182 -16 186 -12
rect 113 -28 114 -26
rect 116 -28 117 -26
rect 113 -30 117 -28
rect 120 -20 136 -19
rect 120 -22 132 -20
rect 134 -22 136 -20
rect 182 -18 183 -16
rect 185 -18 186 -16
rect 182 -20 186 -18
rect 120 -23 136 -22
rect 120 -34 124 -23
rect 110 -35 124 -34
rect 110 -37 112 -35
rect 114 -37 124 -35
rect 110 -38 124 -37
rect 127 -29 131 -27
rect 127 -31 128 -29
rect 130 -31 131 -29
rect 127 -34 131 -31
rect 127 -38 138 -34
rect 120 -42 124 -38
rect 103 -46 112 -42
rect 120 -46 130 -42
rect 54 -54 83 -50
rect 97 -50 103 -49
rect 97 -52 99 -50
rect 101 -52 103 -50
rect 78 -56 79 -54
rect 81 -56 82 -54
rect 78 -58 82 -56
rect 46 -60 56 -59
rect 46 -62 52 -60
rect 54 -62 56 -60
rect 46 -63 56 -62
rect 68 -60 72 -58
rect 68 -62 69 -60
rect 71 -62 72 -60
rect 68 -68 72 -62
rect 97 -68 103 -52
rect 108 -50 112 -46
rect 108 -52 109 -50
rect 111 -51 122 -50
rect 111 -52 118 -51
rect 108 -53 118 -52
rect 120 -53 122 -51
rect 108 -54 122 -53
rect 114 -60 118 -58
rect 114 -62 115 -60
rect 117 -62 118 -60
rect 114 -68 118 -62
rect 126 -59 130 -46
rect 134 -45 138 -38
rect 134 -47 135 -45
rect 137 -47 138 -45
rect 158 -24 163 -22
rect 158 -26 159 -24
rect 161 -26 163 -24
rect 158 -28 163 -26
rect 134 -50 138 -47
rect 159 -50 163 -28
rect 186 -26 190 -24
rect 186 -28 187 -26
rect 189 -28 190 -26
rect 186 -42 190 -28
rect 196 -26 200 -12
rect 262 -16 266 -12
rect 196 -28 197 -26
rect 199 -28 200 -26
rect 196 -30 200 -28
rect 203 -20 219 -19
rect 203 -22 215 -20
rect 217 -22 219 -20
rect 262 -18 263 -16
rect 265 -18 266 -16
rect 262 -20 266 -18
rect 203 -23 219 -22
rect 203 -34 207 -23
rect 193 -35 207 -34
rect 193 -37 195 -35
rect 197 -37 207 -35
rect 193 -38 207 -37
rect 210 -29 214 -27
rect 210 -31 211 -29
rect 213 -31 214 -29
rect 210 -34 214 -31
rect 210 -38 221 -34
rect 203 -42 207 -38
rect 186 -46 195 -42
rect 203 -46 213 -42
rect 134 -54 163 -50
rect 180 -50 186 -49
rect 180 -52 182 -50
rect 184 -52 186 -50
rect 158 -56 159 -54
rect 161 -56 162 -54
rect 158 -58 162 -56
rect 126 -60 136 -59
rect 126 -62 132 -60
rect 134 -62 136 -60
rect 126 -63 136 -62
rect 148 -60 152 -58
rect 148 -62 149 -60
rect 151 -62 152 -60
rect 148 -68 152 -62
rect 180 -68 186 -52
rect 191 -50 195 -46
rect 191 -52 192 -50
rect 194 -51 205 -50
rect 194 -52 201 -51
rect 191 -53 201 -52
rect 203 -53 205 -51
rect 191 -54 205 -53
rect 197 -60 201 -58
rect 197 -62 198 -60
rect 200 -62 201 -60
rect 197 -68 201 -62
rect 209 -59 213 -46
rect 217 -45 221 -38
rect 217 -47 218 -45
rect 220 -47 221 -45
rect 241 -24 246 -22
rect 241 -26 242 -24
rect 244 -26 246 -24
rect 241 -28 246 -26
rect 217 -50 221 -47
rect 242 -50 246 -28
rect 266 -26 270 -24
rect 266 -28 267 -26
rect 269 -28 270 -26
rect 266 -42 270 -28
rect 276 -26 280 -12
rect 276 -28 277 -26
rect 279 -28 280 -26
rect 276 -30 280 -28
rect 283 -20 299 -19
rect 283 -22 295 -20
rect 297 -22 299 -20
rect 283 -23 299 -22
rect 283 -34 287 -23
rect 273 -35 287 -34
rect 273 -37 275 -35
rect 277 -37 287 -35
rect 273 -38 287 -37
rect 290 -29 294 -27
rect 290 -31 291 -29
rect 293 -31 294 -29
rect 290 -34 294 -31
rect 290 -38 301 -34
rect 283 -42 287 -38
rect 266 -46 275 -42
rect 283 -46 293 -42
rect 217 -54 246 -50
rect 260 -50 266 -49
rect 260 -52 262 -50
rect 264 -52 266 -50
rect 241 -56 242 -54
rect 244 -56 245 -54
rect 241 -58 245 -56
rect 209 -60 219 -59
rect 209 -62 215 -60
rect 217 -62 219 -60
rect 209 -63 219 -62
rect 231 -60 235 -58
rect 231 -62 232 -60
rect 234 -62 235 -60
rect 231 -68 235 -62
rect 260 -68 266 -52
rect 271 -50 275 -46
rect 271 -52 272 -50
rect 274 -51 285 -50
rect 274 -52 281 -51
rect 271 -53 281 -52
rect 283 -53 285 -51
rect 271 -54 285 -53
rect 277 -60 281 -58
rect 277 -62 278 -60
rect 280 -62 281 -60
rect 277 -68 281 -62
rect 289 -59 293 -46
rect 297 -45 301 -38
rect 297 -47 298 -45
rect 300 -47 301 -45
rect 321 -24 326 -22
rect 321 -26 322 -24
rect 324 -26 326 -24
rect 321 -28 326 -26
rect 297 -50 301 -47
rect 322 -50 326 -28
rect 297 -54 326 -50
rect 321 -56 322 -54
rect 324 -56 325 -54
rect 321 -58 325 -56
rect 289 -60 299 -59
rect 289 -62 295 -60
rect 297 -62 299 -60
rect 289 -63 299 -62
rect 311 -60 315 -58
rect 311 -62 312 -60
rect 314 -62 315 -60
rect 311 -68 315 -62
rect -61 -115 -60 -109
rect -57 -110 -53 -89
rect -34 -107 -30 -89
rect -34 -109 -33 -107
rect -31 -109 -30 -107
rect -57 -111 -49 -110
rect -57 -113 -53 -111
rect -51 -113 -49 -111
rect -57 -114 -49 -113
rect -45 -111 -39 -110
rect -34 -111 -30 -109
rect -45 -113 -43 -111
rect -41 -113 -39 -111
rect -45 -119 -39 -113
rect -58 -120 -39 -119
rect -58 -122 -56 -120
rect -54 -122 -39 -120
rect -58 -123 -39 -122
rect -61 -134 -60 -132
rect -49 -136 -45 -123
rect -49 -137 -30 -136
rect -49 -139 -34 -137
rect -32 -139 -30 -137
rect -49 -140 -30 -139
rect -49 -177 -30 -176
rect -49 -179 -34 -177
rect -32 -179 -30 -177
rect -49 -180 -30 -179
rect -61 -184 -60 -182
rect -49 -193 -45 -180
rect -58 -194 -39 -193
rect -58 -196 -56 -194
rect -54 -196 -39 -194
rect -58 -197 -39 -196
rect -61 -207 -60 -201
rect -57 -203 -49 -202
rect -57 -205 -53 -203
rect -51 -205 -49 -203
rect -57 -206 -49 -205
rect -45 -203 -39 -197
rect -45 -205 -43 -203
rect -41 -205 -39 -203
rect -45 -206 -39 -205
rect -57 -227 -53 -206
rect -34 -207 -30 -205
rect -34 -209 -33 -207
rect -31 -209 -30 -207
rect -34 -227 -30 -209
rect 17 -110 23 -94
rect 34 -100 38 -94
rect 34 -102 35 -100
rect 37 -102 38 -100
rect 34 -104 38 -102
rect 46 -100 56 -99
rect 46 -102 52 -100
rect 54 -102 56 -100
rect 46 -103 56 -102
rect 68 -100 72 -94
rect 68 -102 69 -100
rect 71 -102 72 -100
rect 17 -112 19 -110
rect 21 -112 23 -110
rect 17 -113 23 -112
rect 28 -109 42 -108
rect 28 -110 38 -109
rect 28 -112 29 -110
rect 31 -111 38 -110
rect 40 -111 42 -109
rect 31 -112 42 -111
rect 28 -116 32 -112
rect 46 -116 50 -103
rect 68 -104 72 -102
rect 78 -106 82 -104
rect 78 -108 79 -106
rect 81 -108 82 -106
rect 23 -120 32 -116
rect 40 -120 50 -116
rect 54 -112 83 -108
rect 54 -115 58 -112
rect 54 -117 55 -115
rect 57 -117 58 -115
rect 23 -134 27 -120
rect 40 -124 44 -120
rect 54 -124 58 -117
rect 30 -125 44 -124
rect 30 -127 32 -125
rect 34 -127 44 -125
rect 30 -128 44 -127
rect 23 -136 24 -134
rect 26 -136 27 -134
rect 23 -138 27 -136
rect 33 -134 37 -132
rect 33 -136 34 -134
rect 36 -136 37 -134
rect 19 -144 23 -142
rect 19 -146 20 -144
rect 22 -146 23 -144
rect 19 -150 23 -146
rect 33 -150 37 -136
rect 40 -139 44 -128
rect 47 -128 58 -124
rect 47 -131 51 -128
rect 47 -133 48 -131
rect 50 -133 51 -131
rect 47 -135 51 -133
rect 40 -140 56 -139
rect 79 -134 83 -112
rect 97 -110 103 -94
rect 114 -100 118 -94
rect 114 -102 115 -100
rect 117 -102 118 -100
rect 114 -104 118 -102
rect 126 -100 136 -99
rect 126 -102 132 -100
rect 134 -102 136 -100
rect 126 -103 136 -102
rect 148 -100 152 -94
rect 148 -102 149 -100
rect 151 -102 152 -100
rect 97 -112 99 -110
rect 101 -112 103 -110
rect 97 -113 103 -112
rect 108 -109 122 -108
rect 108 -110 118 -109
rect 108 -112 109 -110
rect 111 -111 118 -110
rect 120 -111 122 -109
rect 111 -112 122 -111
rect 78 -136 83 -134
rect 78 -138 79 -136
rect 81 -138 83 -136
rect 78 -140 83 -138
rect 108 -116 112 -112
rect 126 -116 130 -103
rect 148 -104 152 -102
rect 158 -106 162 -104
rect 158 -108 159 -106
rect 161 -108 162 -106
rect 103 -120 112 -116
rect 120 -120 130 -116
rect 134 -112 163 -108
rect 134 -115 138 -112
rect 134 -117 135 -115
rect 137 -117 138 -115
rect 103 -134 107 -120
rect 120 -124 124 -120
rect 134 -124 138 -117
rect 110 -125 124 -124
rect 110 -127 112 -125
rect 114 -127 124 -125
rect 110 -128 124 -127
rect 103 -136 104 -134
rect 106 -136 107 -134
rect 40 -142 52 -140
rect 54 -142 56 -140
rect 40 -143 56 -142
rect 103 -138 107 -136
rect 113 -134 117 -132
rect 113 -136 114 -134
rect 116 -136 117 -134
rect 99 -144 103 -142
rect 99 -146 100 -144
rect 102 -146 103 -144
rect 99 -150 103 -146
rect 113 -150 117 -136
rect 120 -139 124 -128
rect 127 -128 138 -124
rect 127 -131 131 -128
rect 127 -133 128 -131
rect 130 -133 131 -131
rect 127 -135 131 -133
rect 120 -140 136 -139
rect 159 -134 163 -112
rect 177 -110 183 -94
rect 194 -100 198 -94
rect 194 -102 195 -100
rect 197 -102 198 -100
rect 194 -104 198 -102
rect 206 -100 216 -99
rect 206 -102 212 -100
rect 214 -102 216 -100
rect 206 -103 216 -102
rect 228 -100 232 -94
rect 228 -102 229 -100
rect 231 -102 232 -100
rect 177 -112 179 -110
rect 181 -112 183 -110
rect 177 -113 183 -112
rect 188 -109 202 -108
rect 188 -110 198 -109
rect 188 -112 189 -110
rect 191 -111 198 -110
rect 200 -111 202 -109
rect 191 -112 202 -111
rect 158 -136 163 -134
rect 158 -138 159 -136
rect 161 -138 163 -136
rect 158 -140 163 -138
rect 188 -116 192 -112
rect 206 -116 210 -103
rect 228 -104 232 -102
rect 238 -106 242 -104
rect 238 -108 239 -106
rect 241 -108 242 -106
rect 183 -120 192 -116
rect 200 -120 210 -116
rect 214 -112 243 -108
rect 214 -115 218 -112
rect 214 -117 215 -115
rect 217 -117 218 -115
rect 183 -134 187 -120
rect 200 -124 204 -120
rect 214 -124 218 -117
rect 190 -125 204 -124
rect 190 -127 192 -125
rect 194 -127 204 -125
rect 190 -128 204 -127
rect 183 -136 184 -134
rect 186 -136 187 -134
rect 120 -142 132 -140
rect 134 -142 136 -140
rect 120 -143 136 -142
rect 183 -138 187 -136
rect 193 -134 197 -132
rect 193 -136 194 -134
rect 196 -136 197 -134
rect 179 -144 183 -142
rect 179 -146 180 -144
rect 182 -146 183 -144
rect 179 -150 183 -146
rect 193 -150 197 -136
rect 200 -139 204 -128
rect 207 -128 218 -124
rect 207 -131 211 -128
rect 207 -133 208 -131
rect 210 -133 211 -131
rect 207 -135 211 -133
rect 200 -140 216 -139
rect 239 -134 243 -112
rect 257 -110 263 -94
rect 274 -100 278 -94
rect 274 -102 275 -100
rect 277 -102 278 -100
rect 274 -104 278 -102
rect 286 -100 296 -99
rect 286 -102 292 -100
rect 294 -102 296 -100
rect 286 -103 296 -102
rect 308 -100 312 -94
rect 308 -102 309 -100
rect 311 -102 312 -100
rect 257 -112 259 -110
rect 261 -112 263 -110
rect 257 -113 263 -112
rect 268 -109 282 -108
rect 268 -110 278 -109
rect 268 -112 269 -110
rect 271 -111 278 -110
rect 280 -111 282 -109
rect 271 -112 282 -111
rect 238 -136 243 -134
rect 238 -138 239 -136
rect 241 -138 243 -136
rect 238 -140 243 -138
rect 268 -116 272 -112
rect 286 -116 290 -103
rect 308 -104 312 -102
rect 318 -106 322 -104
rect 318 -108 319 -106
rect 321 -108 322 -106
rect 263 -120 272 -116
rect 280 -120 290 -116
rect 294 -112 323 -108
rect 294 -115 298 -112
rect 294 -117 295 -115
rect 297 -117 298 -115
rect 263 -134 267 -120
rect 280 -124 284 -120
rect 294 -124 298 -117
rect 270 -125 284 -124
rect 270 -127 272 -125
rect 274 -127 284 -125
rect 270 -128 284 -127
rect 263 -136 264 -134
rect 266 -136 267 -134
rect 200 -142 212 -140
rect 214 -142 216 -140
rect 200 -143 216 -142
rect 263 -138 267 -136
rect 273 -134 277 -132
rect 273 -136 274 -134
rect 276 -136 277 -134
rect 259 -144 263 -142
rect 259 -146 260 -144
rect 262 -146 263 -144
rect 259 -150 263 -146
rect 273 -150 277 -136
rect 280 -139 284 -128
rect 287 -128 298 -124
rect 287 -131 291 -128
rect 287 -133 288 -131
rect 290 -133 291 -131
rect 287 -135 291 -133
rect 280 -140 296 -139
rect 319 -134 323 -112
rect 318 -136 323 -134
rect 318 -138 319 -136
rect 321 -138 323 -136
rect 318 -140 323 -138
rect 280 -142 292 -140
rect 294 -142 296 -140
rect 280 -143 296 -142
rect 19 -176 23 -172
rect 19 -178 20 -176
rect 22 -178 23 -176
rect 19 -180 23 -178
rect 23 -186 27 -184
rect 23 -188 24 -186
rect 26 -188 27 -186
rect 23 -202 27 -188
rect 33 -186 37 -172
rect 99 -176 103 -172
rect 33 -188 34 -186
rect 36 -188 37 -186
rect 33 -190 37 -188
rect 40 -180 56 -179
rect 40 -182 52 -180
rect 54 -182 56 -180
rect 99 -178 100 -176
rect 102 -178 103 -176
rect 99 -180 103 -178
rect 40 -183 56 -182
rect 40 -194 44 -183
rect 30 -195 44 -194
rect 30 -197 32 -195
rect 34 -197 44 -195
rect 30 -198 44 -197
rect 47 -189 51 -187
rect 47 -191 48 -189
rect 50 -191 51 -189
rect 47 -194 51 -191
rect 47 -198 58 -194
rect 40 -202 44 -198
rect 23 -206 32 -202
rect 40 -206 50 -202
rect 17 -210 23 -209
rect 17 -212 19 -210
rect 21 -212 23 -210
rect 17 -228 23 -212
rect 28 -210 32 -206
rect 28 -212 29 -210
rect 31 -211 42 -210
rect 31 -212 38 -211
rect 28 -213 38 -212
rect 40 -213 42 -211
rect 28 -214 42 -213
rect 34 -220 38 -218
rect 34 -222 35 -220
rect 37 -222 38 -220
rect 34 -228 38 -222
rect 46 -219 50 -206
rect 54 -205 58 -198
rect 54 -207 55 -205
rect 57 -207 58 -205
rect 78 -184 83 -182
rect 78 -186 79 -184
rect 81 -186 83 -184
rect 78 -188 83 -186
rect 54 -210 58 -207
rect 79 -210 83 -188
rect 103 -186 107 -184
rect 103 -188 104 -186
rect 106 -188 107 -186
rect 103 -202 107 -188
rect 113 -186 117 -172
rect 179 -176 183 -172
rect 113 -188 114 -186
rect 116 -188 117 -186
rect 113 -190 117 -188
rect 120 -180 136 -179
rect 120 -182 132 -180
rect 134 -182 136 -180
rect 179 -178 180 -176
rect 182 -178 183 -176
rect 179 -180 183 -178
rect 120 -183 136 -182
rect 120 -194 124 -183
rect 110 -195 124 -194
rect 110 -197 112 -195
rect 114 -197 124 -195
rect 110 -198 124 -197
rect 127 -189 131 -187
rect 127 -191 128 -189
rect 130 -191 131 -189
rect 127 -194 131 -191
rect 127 -198 138 -194
rect 120 -202 124 -198
rect 103 -206 112 -202
rect 120 -206 130 -202
rect 54 -214 83 -210
rect 97 -210 103 -209
rect 97 -212 99 -210
rect 101 -212 103 -210
rect 78 -216 79 -214
rect 81 -216 82 -214
rect 78 -218 82 -216
rect 46 -220 56 -219
rect 46 -222 52 -220
rect 54 -222 56 -220
rect 46 -223 56 -222
rect 68 -220 72 -218
rect 68 -222 69 -220
rect 71 -222 72 -220
rect 68 -228 72 -222
rect 97 -228 103 -212
rect 108 -210 112 -206
rect 108 -212 109 -210
rect 111 -211 122 -210
rect 111 -212 118 -211
rect 108 -213 118 -212
rect 120 -213 122 -211
rect 108 -214 122 -213
rect 114 -220 118 -218
rect 114 -222 115 -220
rect 117 -222 118 -220
rect 114 -228 118 -222
rect 126 -219 130 -206
rect 134 -205 138 -198
rect 134 -207 135 -205
rect 137 -207 138 -205
rect 158 -184 163 -182
rect 158 -186 159 -184
rect 161 -186 163 -184
rect 158 -188 163 -186
rect 134 -210 138 -207
rect 159 -210 163 -188
rect 183 -186 187 -184
rect 183 -188 184 -186
rect 186 -188 187 -186
rect 183 -202 187 -188
rect 193 -186 197 -172
rect 259 -176 263 -172
rect 193 -188 194 -186
rect 196 -188 197 -186
rect 193 -190 197 -188
rect 200 -180 216 -179
rect 200 -182 212 -180
rect 214 -182 216 -180
rect 259 -178 260 -176
rect 262 -178 263 -176
rect 259 -180 263 -178
rect 200 -183 216 -182
rect 200 -194 204 -183
rect 190 -195 204 -194
rect 190 -197 192 -195
rect 194 -197 204 -195
rect 190 -198 204 -197
rect 207 -189 211 -187
rect 207 -191 208 -189
rect 210 -191 211 -189
rect 207 -194 211 -191
rect 207 -198 218 -194
rect 200 -202 204 -198
rect 183 -206 192 -202
rect 200 -206 210 -202
rect 134 -214 163 -210
rect 177 -210 183 -209
rect 177 -212 179 -210
rect 181 -212 183 -210
rect 158 -216 159 -214
rect 161 -216 162 -214
rect 158 -218 162 -216
rect 126 -220 136 -219
rect 126 -222 132 -220
rect 134 -222 136 -220
rect 126 -223 136 -222
rect 148 -220 152 -218
rect 148 -222 149 -220
rect 151 -222 152 -220
rect 148 -228 152 -222
rect 177 -228 183 -212
rect 188 -210 192 -206
rect 188 -212 189 -210
rect 191 -211 202 -210
rect 191 -212 198 -211
rect 188 -213 198 -212
rect 200 -213 202 -211
rect 188 -214 202 -213
rect 194 -220 198 -218
rect 194 -222 195 -220
rect 197 -222 198 -220
rect 194 -228 198 -222
rect 206 -219 210 -206
rect 214 -205 218 -198
rect 214 -207 215 -205
rect 217 -207 218 -205
rect 238 -184 243 -182
rect 238 -186 239 -184
rect 241 -186 243 -184
rect 238 -188 243 -186
rect 214 -210 218 -207
rect 239 -210 243 -188
rect 263 -186 267 -184
rect 263 -188 264 -186
rect 266 -188 267 -186
rect 263 -202 267 -188
rect 273 -186 277 -172
rect 273 -188 274 -186
rect 276 -188 277 -186
rect 273 -190 277 -188
rect 280 -180 296 -179
rect 280 -182 292 -180
rect 294 -182 296 -180
rect 280 -183 296 -182
rect 280 -194 284 -183
rect 270 -195 284 -194
rect 270 -197 272 -195
rect 274 -197 284 -195
rect 270 -198 284 -197
rect 287 -189 291 -187
rect 287 -191 288 -189
rect 290 -191 291 -189
rect 287 -194 291 -191
rect 287 -198 298 -194
rect 280 -202 284 -198
rect 263 -206 272 -202
rect 280 -206 290 -202
rect 214 -214 243 -210
rect 257 -210 263 -209
rect 257 -212 259 -210
rect 261 -212 263 -210
rect 238 -216 239 -214
rect 241 -216 242 -214
rect 238 -218 242 -216
rect 206 -220 216 -219
rect 206 -222 212 -220
rect 214 -222 216 -220
rect 206 -223 216 -222
rect 228 -220 232 -218
rect 228 -222 229 -220
rect 231 -222 232 -220
rect 228 -228 232 -222
rect 257 -228 263 -212
rect 268 -210 272 -206
rect 268 -212 269 -210
rect 271 -211 282 -210
rect 271 -212 278 -211
rect 268 -213 278 -212
rect 280 -213 282 -211
rect 268 -214 282 -213
rect 274 -220 278 -218
rect 274 -222 275 -220
rect 277 -222 278 -220
rect 274 -228 278 -222
rect 286 -219 290 -206
rect 294 -205 298 -198
rect 294 -207 295 -205
rect 297 -207 298 -205
rect 318 -184 323 -182
rect 318 -186 319 -184
rect 321 -186 323 -184
rect 318 -188 323 -186
rect 294 -210 298 -207
rect 319 -210 323 -188
rect 294 -214 323 -210
rect 318 -216 319 -214
rect 321 -216 322 -214
rect 318 -218 322 -216
rect 286 -220 296 -219
rect 286 -222 292 -220
rect 294 -222 296 -220
rect 286 -223 296 -222
rect 308 -220 312 -218
rect 308 -222 309 -220
rect 311 -222 312 -220
rect 308 -228 312 -222
<< via1 >>
rect -101 35 -99 37
rect -66 36 -64 38
rect -80 27 -78 29
rect -91 7 -89 9
rect -92 -20 -90 -18
rect -39 28 -37 30
rect -29 8 -27 10
rect -70 -5 -68 -3
rect -80 -27 -78 -25
rect -38 -27 -36 -25
rect -65 -36 -63 -34
rect -47 -59 -45 -57
rect 72 34 74 36
rect 154 34 156 36
rect 235 34 237 36
rect 318 34 320 36
rect 4 8 6 10
rect 72 -35 74 -33
rect 152 -35 154 -33
rect 235 -35 237 -33
rect 315 -35 317 -33
rect -151 -131 -149 -129
rect -46 -98 -44 -96
rect -64 -121 -62 -119
rect -37 -130 -35 -128
rect -27 -167 -25 -165
rect -151 -188 -149 -186
rect -37 -188 -35 -186
rect -64 -211 -62 -209
rect -163 -221 -161 -219
rect -46 -220 -44 -218
rect 72 -129 74 -127
rect 152 -129 154 -127
rect 232 -129 234 -127
rect 312 -129 314 -127
rect 4 -167 6 -165
rect 72 -195 74 -193
rect 152 -195 154 -193
rect 232 -195 234 -193
rect 312 -195 314 -193
<< labels >>
rlabel alu1 191 70 196 76 0 vdd
rlabel alu1 28 -75 33 -69 0 vdd
rlabel alu1 190 -75 195 -69 0 vdd
rlabel alu1 29 -93 34 -87 0 vdd
rlabel alu1 190 -93 195 -87 0 vdd
rlabel alu1 26 -235 31 -229 0 vdd
rlabel alu1 267 -235 272 -229 0 vdd
rlabel alu1 39 -171 44 -165 0 vss
rlabel alu1 162 -171 167 -165 0 vss
rlabel alu1 41 -157 46 -151 0 vss
rlabel alu1 241 -157 246 -151 0 vss
rlabel alu1 45 -11 50 -5 0 vss
rlabel alu1 215 -11 220 -5 0 vss
rlabel alu1 46 6 51 12 0 vss
rlabel alu1 216 6 221 12 0 vss
rlabel alu1 82 70 87 76 0 vdd
rlabel nwell -123 67 -116 75 0 vdd
rlabel alu1 -124 -76 -117 -68 0 vdd
rlabel nwell -52 70 -45 78 0 vdd
rlabel nwell -52 -74 -45 -66 0 vdd
rlabel nwell -52 -89 -45 -81 0 vdd
rlabel nwell -52 -235 -45 -227 0 vdd
rlabel pwell -123 3 -116 11 0 vss
rlabel pwell -124 -12 -117 -4 0 vss
rlabel alu1 -36 5 -29 13 0 vss
rlabel alu1 -35 -10 -28 -2 0 vss
rlabel alu1 -36 -153 -29 -145 0 vss
rlabel alu1 -35 -171 -28 -163 0 vss
rlabel space -146 56 -139 64 0 a
rlabel space -148 -63 -141 -55 0 b
rlabel alu2 -49 -59 -49 -59 1 a
rlabel alu2 -47 -220 -47 -220 1 a
rlabel alu2 -39 -130 -39 -130 1 b
rlabel alu2 -38 -186 -38 -186 1 b
rlabel alu1 -127 34 -127 34 1 inv1
rlabel alu1 -50 61 -50 61 1 inv1
rlabel alu2 -48 -99 -48 -99 1 inv1
rlabel alu1 -126 -36 -126 -36 1 inv2
rlabel alu2 -42 28 -42 28 1 inv2
rlabel alu2 -41 -26 -41 -26 1 inv2
rlabel pdifct1 -65 45 -65 45 1 D0
rlabel alu1 -64 -45 -64 -45 1 D1
rlabel alu1 -63 -115 -63 -115 1 D2
rlabel alu1 -63 -193 -63 -193 1 D3
rlabel alu1 73 25 73 25 1 D0
rlabel alu1 155 24 155 24 1 D0
rlabel alu1 236 22 236 22 1 D0
rlabel alu1 319 23 319 23 1 D0
rlabel alu1 63 29 63 29 1 R03
rlabel alu1 9 27 9 27 1 O03
rlabel alu1 92 28 92 28 1 O02
rlabel alu1 144 29 144 29 1 R02
rlabel alu1 224 29 224 29 1 R01
rlabel alu1 173 28 173 28 1 O01
rlabel alu1 307 29 307 29 1 R00
rlabel alu1 256 28 256 28 1 O00
rlabel alu1 73 -21 73 -21 1 D1
rlabel alu1 62 -28 62 -28 1 R13
rlabel alu1 9 -28 9 -28 1 O13
rlabel alu1 152 -21 152 -21 1 D1
rlabel alu1 141 -29 141 -29 1 R12
rlabel alu1 90 -28 90 -28 1 O12
rlabel alu1 235 -22 235 -22 1 D1
rlabel alu1 224 -28 224 -28 1 R11
rlabel alu1 173 -28 173 -28 1 O11
rlabel alu1 315 -20 315 -20 1 D1
rlabel alu1 303 -28 303 -28 1 R10
rlabel alu1 253 -27 253 -27 1 O10
rlabel alu1 73 -138 73 -138 1 D2
rlabel alu1 61 -134 61 -134 1 R23
rlabel alu1 10 -134 10 -134 1 O23
rlabel alu1 153 -142 153 -142 1 D2
rlabel alu1 141 -134 141 -134 1 R22
rlabel alu1 90 -134 90 -134 1 O22
rlabel alu1 233 -141 233 -141 1 D2
rlabel alu1 221 -134 221 -134 1 R21
rlabel alu1 169 -135 169 -135 1 O21
rlabel alu1 313 -141 313 -141 1 D2
rlabel alu1 302 -134 302 -134 1 R20
rlabel alu1 250 -134 250 -134 1 O20
rlabel alu1 73 -181 73 -181 1 D3
rlabel alu1 61 -188 61 -188 1 R33
rlabel alu1 10 -187 10 -187 1 O33
rlabel alu1 152 -181 152 -181 1 D3
rlabel alu1 141 -188 141 -188 1 R32
rlabel alu1 89 -188 89 -188 1 O32
rlabel alu1 233 -181 233 -181 1 D3
rlabel alu1 221 -188 221 -188 1 R31
rlabel alu1 170 -186 170 -186 1 R30
rlabel alu1 313 -181 313 -181 1 D3
rlabel alu1 302 -188 302 -188 1 R30
rlabel alu1 250 -188 250 -188 1 O30
<< end >>
