* ===============================
* 1-Word x 4-Bit ROM Demo
* Using active-high 2-to-4 decoder
* ===============================

* --- Power Supply ---
Vdd vdd 0 5

* --- Address Inputs ---
Va a 0 PULSE(0 5 0 5n 5n 20n 40n)   ; MSB
Vb b 0 PULSE(0 5 0 5n 5n 40n 80n)   ; LSB

* --- Include transistor models ---
.include "t14y_tsmc_025_level3.txt"

* ===============================
* 2-to-4 Decoder Subcircuit
* ===============================
.subckt DEC2to4 A B Y0 Y1 Y2 Y3 vdd gnd

* --- Inverters for Abar and Bbar ---
Mp1 Abar A vdd vdd CMOSP W=4u L=1u
Mn1 Abar A 0   0   CMOSN W=2u L=1u
Mp2 Bbar B vdd vdd CMOSP W=4u L=1u
Mn2 Bbar B 0   0   CMOSN W=2u L=1u

* --- NAND-style outputs (active-low) ---
* Y0 = Abar & Bbar
Mp3 Y0 Abar vdd vdd CMOSP W=4u L=1u
Mp4 Y0 Bbar vdd vdd CMOSP W=4u L=1u
Mn3 Y0 Abar n1 n1 CMOSN W=2u L=1u
Mn4 n1 Bbar 0   0   CMOSN W=2u L=1u

* Y1 = Abar & B
Mp5 Y1 Abar vdd vdd CMOSP W=4u L=1u
Mp6 Y1 B    vdd vdd CMOSP W=4u L=1u
Mn5 Y1 Abar n2 n2 CMOSN W=2u L=1u
Mn6 n2 B    0   0  CMOSN W=2u L=1u

* Y2 = A & Bbar
Mp7 Y2 A vdd vdd CMOSP W=4u L=1u
Mp8 Y2 Bbar vdd vdd CMOSP W=4u L=1u
Mn7 Y2 A n3 n3 CMOSN W=2u L=1u
Mn8 n3 Bbar 0   0  CMOSN W=2u L=1u

* Y3 = A & B
Mp9  Y3 A vdd vdd CMOSP W=4u L=1u
Mp10 Y3 B vdd vdd CMOSP W=4u L=1u
Mn9  Y3 A n4 n4 CMOSN W=2u L=1u
Mn10 n4 B 0   0 CMOSN W=2u L=1u

* --- Active-High Outputs (wordlines) ---
Myn0 Y0h Y0 0 0 CMOSN W=2u L=1u
Myp0 Y0h Y0 vdd vdd CMOSP W=4u L=1u

Myn1 Y1h Y1 0 0 CMOSN W=2u L=1u
Myp1 Y1h Y1 vdd vdd CMOSP W=4u L=1u

Myn2 Y2h Y2 0 0 CMOSN W=2u L=1u
Myp2 Y2h Y2 vdd vdd CMOSP W=4u L=1u

Myn3 Y3h Y3 0 0 CMOSN W=2u L=1u
Myp3 Y3h Y3 vdd vdd CMOSP W=4u L=1u

.ends DEC2to4

* ===============================
* Instantiate Decoder
* ===============================
Xdec a b Y0 Y1 Y2 Y3 vdd 0 DEC2to4

* ===============================
* Single ROM Word (1 row, 4 bits)
* Stored Data: 1 0 1 1 (example)
* ===============================

* ROM cells connected to active-high wordline Y0h
* Pass transistor connecting stored value to bitline when wordline = 1
* Bit0 = 1
Mcell0 BL0 vdd Y0h 0 CMOSN W=2u L=1u
* Bit1 = 0
Mcell1 BL1 0   Y0h 0 CMOSN W=2u L=1u
* Bit2 = 1
Mcell2 BL2 vdd Y0h 0 CMOSN W=2u L=1u
* Bit3 = 1
Mcell3 BL3 vdd Y0h 0 CMOSN W=2u L=1u

* Output Buffers (optional, strengthens bitline signals)
Mbuf0_out OUT0 BL0 0 0 CMOSN W=2u L=1u
Mbuf0_p   OUT0 BL0 vdd vdd CMOSP W=4u L=1u

Mbuf1_out OUT1 BL1 0 0 CMOSN W=2u L=1u
Mbuf1_p   OUT1 BL1 vdd vdd CMOSP W=4u L=1u

Mbuf2_out OUT2 BL2 0 0 CMOSN W=2u L=1u
Mbuf2_p   OUT2 BL2 vdd vdd CMOSP W=4u L=1u

Mbuf3_out OUT3 BL3 0 0 CMOSN W=2u L=1u
Mbuf3_p   OUT3 BL3 vdd vdd CMOSP W=4u L=1u

* ===============================
* Simulation
* ===============================
.tran 1n 200n
.probe v(a) v(b) v(Y0h) v(OUT0) v(OUT1) v(OUT2) v(OUT3)
plot v(a) v(b) v(Y0h) v(OUT0) v(OUT1) v(OUT2) v(OUT3)
.end
