* 1-Word x 4-Bit ROM Demo

* --- Power Supply ---
Vdd vdd 0 5

* --- Address Inputs ---
Va a 0 PULSE(0 5 0 5n 5n 20n 40n)
Vb b 0 PULSE(0 5 0 5n 5n 40n 80n)

* --- Include transistor models ---
.include "t14y_tsmc_025_level3.txt"

* --- Include decoder subcircuit ---
.include "DEC2to4.cir"

* --- Instantiate decoder ---
Xdec a b Y0 Y1 Y2 Y3 vdd 0 DEC2to4

* --- ROM Cells (1 Word x 4 bits example) ---
Mcell0 BL0 vdd Y0h 0 CMOSN W=2u L=1u   ; Bit0=1
Mcell1 BL1 0   Y0h 0 CMOSN W=2u L=1u   ; Bit1=0
Mcell2 BL2 vdd Y0h 0 CMOSN W=2u L=1u   ; Bit2=1
Mcell3 BL3 vdd Y0h 0 CMOSN W=2u L=1u   ; Bit3=1

* --- Output Buffers ---
Mbuf0_out OUT0 BL0 0 0 CMOSN W=2u L=1u
Mbuf0_p   OUT0 BL0 vdd vdd CMOSP W=4u L=1u
Mbuf1_out OUT1 BL1 0 0 CMOSN W=2u L=1u
Mbuf1_p   OUT1 BL1 vdd vdd CMOSP W=4u L=1u
Mbuf2_out OUT2 BL2 0 0 CMOSN W=2u L=1u
Mbuf2_p   OUT2 BL2 vdd vdd CMOSP W=4u L=1u
Mbuf3_out OUT3 BL3 0 0 CMOSN W=2u L=1u
Mbuf3_p   OUT3 BL3 vdd vdd CMOSP W=4u L=1u

* --- Simulation ---
.tran 1n 200n
.probe v(a) v(b) v(Y0h) v(OUT0) v(OUT1) v(OUT2) v(OUT3)
.end
